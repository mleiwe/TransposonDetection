 tpg|BK006937.2| 316620 + tpg|BK006937.2| 315874 - INS GGTATATACTGTAGCATCCGTGTGCGTATGCCCCATCAATATAAGTGAAGGTGAGTATGGCATGTGGTGGTGGTATAGAGTGGTAGGGTAAGTATGTATGTATTATTTACGATCATTTGTTAACGTTTCAATATGGTGGGTGAACAACAGTACAGTGAGTAGGACATGGTGGATGGTAGGGTAATAGTAGGGTAAGTGGTGGTGGAGTTGGATATGGGTAATTGGAGGGTAACGGTTATGATGGGCGGTGGATGGTGGTAGTAAGTAGAGAGATGGATGGTGGTTGGGAGTGGTATGGTTGAGTGGGGCAGGGTAACGAGTGGGGAGGTAGGGTAATGTGAGGGTAGGTTTGGAGACAGGTAAAATCAGGGTTAGAATAGGGTAGTGTTAGGGTAGTGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGTGGGTGTGGTGGGTGTGGTGTGTGTGTGGGTGTGGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGTGTGTGTGGGTGTGTGGGTGTGTGGGTG tpg|BK006937.2|:314504-316619 7X494=56S 1S1=416S 
 tpg|BK006942.2| 439887 + tpg|BK006942.2| 439256 - INS GTATAGACCGCTGAGGCAAGTACCGTGCACAATGATGTGAGTGCATTTGTACTGATTTAGTGAGAGATGGGCCATGGAGTGGAGTGGAATGTGAGAGTAGGGTAAGTTTGAGAGTGGTATATACTGTAGCATCCGTGTGCGTATGCCCTATCAGTATACAATTAAAGGTGAGTATGGCATGTGGTGGTGGGATTAGAGTGGTAGGGTAAGTATGTGTGTATTATTTACGATCATTTGTTAACGTTTCAATATGGTGGGTAGAACAACAGTATAGTGAGTAGCAGATGGTGGATGGTAGGGTAATGGTAGGGTAAGTGGCAGTGGGGTTGGATATGGGTAATTGGAGGGTAACGGTTATGGTGGACGGTGGGTTGGTGGTAGTACGTAGAGAGATGGATTGTGGTTCGGAGTGGTATGGTTGAATGGAACAGGGTAACAAGTGGGGAGGAAGGGTAATGGAGGGTAAGTTGAGAGACAGGATGGTTAGGGTTAAAGTAGGGTAGTGTTAGGGTAGTGTGGTGTGTGGGTGTGGGTGTGGATGTGGTGTGGATGTGGTGTGGGTGTGGATGTGGGTGTGGTGTGTGTGGGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGGTGTGGGTGTGGTGTGGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGT tpg|BK006942.2|:437658-439887 7X586=107S 5S1=704S 
 tpg|BK006942.2| 333255 + tpg|BK006942.2| 333328 - INS GCCCTAGAGAGTATAAGCGTTTCGTCTCCTCTTCCTTTCTCTACTGCAGATTTTCTTGCTGGTTGTTTGATTTTTTCTTTTTAGTGTTCCCCAGATCCAATTGTTCAACCGCCCACACACAACAATGTCTTTCACTAAAATCGCTGCCTTATTAGCTGTTGCCGCTGCCTCCACTCAATTGGTTTCTGCTGAAGTTGGACAATATGAAATCGTCGAATTTGACGCTATTTTGGCTGATGTCAAGGCCAATTTGGAACAATATATGTCCTTGGCAATGAATAATCCAGACTTTACCCTACCATCTGGTGTTTTGGATGTTTACCAACATATGACCACTGCTACTGATGATTCCTACACCAGTTATTTCACCGAAATGGACTTTGCTCAAATCACCAC tpg|BK006942.2|:332449-334134 7X207= 198=7X 
 tpg|BK006942.2| 257491 + tpg|BK006942.2| 257662 - INS TCTGTACACCGCACTCCTCGGTATCGCAAGTGGAAAAAAGGCAGTAAAGAAGTTTCAATCCTTCAATTCTTTTCAACAGCGATAACTTCCATTTCTAAATCAACATTCAAAGGTAAGGAAGCAACACCAACACAGGATCTTGCAGGCTTATGGGTGTGGAAGTGTTTGGCGTATACAGAGTTGAATTCGGCAAAGTTTTTCATGTCAGCCAAGAATACGTTGACTTTGACTATATTGTCTAAAGAAGAATTACTTTCTGCTAAGATATTCTTAACGTTTTGAAAAACTTGTTCGGCCTTCTCAGAGATAGAACCTTGAACAGGCTTGTTATCTGGAGTATAAGGGATTTGACCAGACACGTACACAAAATTGTTGGCCTTCATAGCTTGGGAGTAAGAGGCGGCAGCGGGTGGGGCCAACTTGGTGC tpg|BK006942.2|:256623-258530 7X4=157S 401=7X 
 tpg|BK006942.2| 344765 + tpg|BK006942.2| 344965 - INS GGTTGATCATGGCTGGTACGAACCAGAATGCAACTGAAATCAGATATACCAGATTCCATTCAACGACGTCTGTTCCCCCTCATTAAAGCAACTTATGCACAAGAGGGACTAAAGGGATTTTATTCTGGATTTACTACTAACCTAGTACGAACCATTCCGGCCTCGGCAATCACTCTAGTGTCCTTTGAGTATTTCAGAAACCGCCTAGAAAATATTAGCACTATGGTAATTTAAAGCCTTAAAATTCACACACGCCACACATTGAGTGTGCTATGAATATGCC tpg|BK006942.2|:344185-345545 7X197= 266=7X 
 tpg|BK006942.2| 188851 + tpg|BK006942.2| 189239 - INS GTTGGATCTATTCCTCACAAAATTGGAGCCACAGTTGCAAAAGCAACTGGAAAATTGTGCATTCCCAATGACTTTGAATTTAGCACTATTGATAACTGCCTGTGAATTTGCGAAGAGAGCATCTAATCATAAAAAATACCGGTATAAAAATACGAGGGATTCCGACATTTGTACTCCAAAGAGTAAGAATACTGCTATCGTTAGCAAATTATCGAATACTAAAACTATAAGTAAGAATAAGGTTATTGAAAAGAGTGATAAGAAAAATTACTTTGATAAGAACAGTCAACACA tpg|BK006942.2|:188251-189839 7X178=41S 1=168S 
 tpg|BK006942.2| 411684 + tpg|BK006942.2| 411731 - INS CTTAACTACAAAGAACATGTGTATGAAATACGTAAGAGTATAAGAGTCTCCCATGTCAAATTAACGATTATTCCAGATGGAGGAGTGAAAAGAATAAGAGTTTGGGGGTACTGATAAATACTTAACTACTGTATATTTTAAACCAATGCACTCTTGGCACTTTAAAAGTAAAGGTATAAATGTAGTTAAAAGTTTTTGTTTTGATAATTGAATGTTTTCATTTCGCTATCCCCACG tpg|BK006942.2|:411198-412217 13S18=445S 118=7X 
 tpg|BK006937.2| 92895 + tpg|BK006937.2| 92480 - INS AAATAAAAAACACTCAATGACCTGACCATTTGATGGAGTTTAAGTCAATACCTTCTTGAACCATTTCCCATAATGGTGAAAGTTCCCTCAAGAATTTTACTCTGTCAGAAACGGCCTTAACGACGTAGTCGATATGGTGCACTCTCAGTACAATCTGCTCTGATGCCGCATAGTTAAGCCAGCCCCGACACCCGCCAACACCCGCTGACGCGCCCTGACGGGCTTGTCTGCTCCCGGCATCCGCTTACAGACAAGCTGTGACCGTCTCCGGGAGCTGCATGTGTCAGAGGTTTTCACCGTCATCACCGAAACGCGCGAGACGAAAGGGCCTCGTGATACGCCTATTTTTATAGGTTAATGTCATGATAATAATGGTTTCTTAGGACGGATCGCTTGCCTGTAACTTACACGCGCCTCGTATCTTTTAATGATGGAATAATTGGGGAATTTACTCTGTGTTTATTTATTTTTATGTTTTGTATTTGGATTTTAGAAAGTAAATAAAGAAGGTAGAAGAGTTACGGAATGAAGAAAAAAAAATAAACAAAGGTTTAAAAAATTTCAACAAAAAGCGTACTTTACATATATAT tpg|BK006937.2|:91286-94089 7X132=163S 443S5=7X 
 tpg|BK006942.2| 75170 + tpg|BK006942.2| 75917 - INS GTTGAAGAAGGAGATGCAGTGGCGGGCGTATTGATTGTGTCGCTAGAGGAATCTAAGGAAAGTAAAGAGGCAAATATGGAGGGCCGCAAACTTAAAGACTTAACTGTTTGGTGTTCGTATGCTGCAGTGACAAAGTATGTCACACAACATCCAAAACTAATTCCTATAGTAATTGAAATGCCCCAAGTGAACC tpg|BK006942.2|:74770-76317 7X2=1X7=86S 92S5=7X 
 tpg|BK006942.2| 288095 + tpg|BK006942.2| 288124 - INS CAAATAGATGAATTATGTTTGCATGACCATTGTGTGGCTGATCAAAGATATAGGGCCTGATGAATTTTAAAACGTCCTCCTTTTGATTTGTGTAATATTGATCTTTTTGAAATGGCAAAGTCGTTGGAGGCACTTTTTCGTTAGACAAATCCGTTAAGATTTTGATTTCTCTCTTGATCTTCTTCTTTTTAACTGGTTTCAACATCTTAATAACAATTTTAACTTTAGAGTCTAATTTGACACCTTGGAAAACCTCGGAGTATTTTCCTCGCCCAACTTTATTTTCAATTTCATAGTCCTTTGTATTTGTGGACCAATCAATTAC tpg|BK006942.2|:287431-288788 7X292=14S 1=337S 
 tpg|BK006942.2| 289607 + tpg|BK006942.2| 289813 - INS CCTCTGACCATACCCTGCATTTCATAGTTCGAATCAAATATTCCTTCTACAACCCCCTATTTTTGTCTGTATATTTGACTTCTTAAGTCCCTATTCAGAAAACTCCTAGTAGGTAATTGCAATACACCGAGTATCAACAGTATATGAAGTCCCTTAATCCGTTTTACTACAGGACTGCGAGGTTCGTCTAATTGCTACTGAAATTTTCCAAGCGTTGGTCATATTTTTGATTTTTCGCTTTTTCTTCAGTGTTCGTTCCGAGTGATTTTTGATAGCGCTTTTCTACCACTTAGTGCTGCTGTATGTATTTATATGATATACCAGCGATACATGTAAATATTTCTATAAA tpg|BK006942.2|:288895-290525 7X236S 328=7X 
 tpg|BK006942.2| 262346 + tpg|BK006942.2| 261691 - INS CATAAAAGTCTTCAAACACAGATACCCATCCTTTGATGTATGATAATCGCCTCTCGCAGGATGATAATTTCAAATTTACTAATATTGCTTCGTCACCACCGTCGTCTTCAAACAATATTTTTTCAAAAGCCCTCTCATATTTAAAAGTATCTAACACAAAAAACTGGTCCAAGTTTGGTTCACCCATAGAACTCAGTGATCAACACATCGAAAGAGAAATACATCCAGACACGACTCCTGTGTACGATAGGAATAGATACGTTTCGAATGAACTATCTAATGCCAAATATAATGCCGTTACTTTTGTGCCAACCCTATTATATGAACAGTTCAAATTCTTTTACAATTTATAC tpg|BK006942.2|:260971-263066 7X5=233S 177=7X 
 tpg|BK006942.2| 339222 + tpg|BK006942.2| 339702 - INS GGCTTGGAGAGCATACATCAAGCCCAATGGAGAACACAAATTCCACATCTTCGCATCTACTTCCCATAAATGGATGAAGATTTTCCTTGGTTGCATATCCCAGGGTATCCCCGTAGTAACCGCGTATGATACTTTGGGTGAGAGCGGTTTGATTCACTCCATGGTTGAAACCGAGTCTGCTGCTATTTTCACTGATAATCAATTATTGGCTAAAATGATAGTGCCTTTGCAATCTGCTAAAG tpg|BK006942.2|:338724-340200 7X6=254S 227=7X 
 tpg|BK006942.2| 438042 + tpg|BK006942.2| 438777 - INS GGAAAGGATAACACGTCATGGTAGTGCTCATACTTCAAGTCAAAGTGTTTATTTCGTAAAGTTGAAAGGTAAAATATTTTTATGTTTAGGTGATTTTAGTGGTAATTTTTCTGTAATATTGACATAAGTTTATAAAAATTGAGTGGTTAGTATATGGCGTAAAAGTGGTATAATGTATGCATTAAGAGCAGTTATACAATATTTGGAGCCGCTGAATGAGATATAGATATTAAAATGTGGATAATCGTGAGCTTTATGGGTAAATGGCACAGGGTATAGAC tpg|BK006942.2|:437466-439353 54S188= 264=7X 
 tpg|BK006942.2| 304104 + tpg|BK006942.2| 304836 - INS GTTGGGTGTTCCTTCAATTTATGTATTTCTCTCCATTTTTCCAGATTCCATGTGGCTAATAACACTAGCATTTTAAAGTTTATTTCTTGAGCGGTACTATCATCAAAATCTTGAAACATTATAGGGATACGGGAAACAAAATTGTTCAAAAACAGTTGCAACAACTCTTCATCAACCTCGATTGGGTAATCCCTGCCAAGAATTGTCAGTTTATTGATGTAGAGCTCGTACAAAGAACAAGTTAAATCTTTGTAGTCGTCCCTAGAATTATTT tpg|BK006942.2|:303544-305396 30S89=24S 128S9=7X 
 tpg|BK006942.2| 204797 + tpg|BK006942.2| 204985 - INS ATTTAGAGCCTATTAGTGTAGGCGTGAGCTCTTATACACAGTTTATGTCGCCTCTACTTTCTTAGCATAATCAGGTTTTTTTCTTGATTTTTTTATCATAAATTGTAACTCCGATTTAAGTAGAAGTGAAAAAAAAAATACCCTGTTAATTGTCACAGCATCACTTCTTCCTGTTACTTTCAAAGCTGTAAAGTGTTAGCA tpg|BK006942.2|:204381-205401 7X8=170S 15S155=7X 
 tpg|BK006942.2| 302750 + tpg|BK006942.2| 302099 - INS CCTTATGGACGATGCAAGGTTATTCAGACGCGTTGTTTGTATGCCATTTCCAATGATAATGTTGGTTGCCTTATATAGAAATGTGTTAGGAAGAGATTCTACAGTTGATTGCAGCTTTGACGTTATACTTACACCTTGGATAATGGCCAGTATGTTTTCCAAACGTATGGTGAATTGGTCTAATCCACGTCAAGCTGTTTTAAAAGTATGCAGCGCAGCCGTGACCTCCCGGATAGTTGCCAATTGGTTGTTTACGATGAACATATTATATACCAGTGGTGAAAAGGGTTTTTACTCGCTAGCAACAGCTGTGGTAATTAAAACGGTCACTGATGGGTTTACGGTGATACGGGTTTTCTCTATTCACCTGAACGAGTCAGTATATAGCAAGCCATTACCATAACATTGGGTAACGTCGCACGCAACACAGCTGCGGGTGTGTGTGGTGATTGGTTAGTCAATTGGTCATTTGGGCTGGTAATAGGG tpg|BK006942.2|:301113-303736 7X5=386S 243=7X 
 tpg|BK006942.2| 421911 + tpg|BK006942.2| 421478 - INS CCTCTTCTTCAAGGGTGCCTCAGACCTGGCTACACCGTAAACAACCGTGTCCTTGTCCAAACTGAAAAGAACATCCACGATGGACTTACCGATACCTCTGGAAACACCTGTAACTAAAATAACTTTACCCATGTTTTTTTAACCTGTTACACGCTGTAGTTAGACCCTTTTTTTTAGGTACAATATTC tpg|BK006942.2|:421088-422301 7X5=211S 94=7X 
 tpg|BK006942.2| 430257 + tpg|BK006942.2| 430952 - INS GAGAAAGTTGTGCCAGAATCCAACATCACTGGAAATTGAATATCCGAAACAGTTTTATTGCCAGATTCACTATCCAAAATTGCCACACTTTGTGCAGTAATAATCATCCCAGGATTTGAGCCAAGGGTATTGAATGCCTGCAGCATAGGCAGGGTGTAAAGC tpg|BK006942.2|:429919-431290 7X81= 181S3=7X 
 tpg|BK006942.2| 138941 + tpg|BK006942.2| 139689 - INS ACTCGACCCTAGGCGCTAGGGTGGGTGACGCATTTTAACTTTGCAACAGAATGCCATATGCGGTGTTAACCTCACAAGATCGGCTCTACTATCTGCAAGCTGCGGCAAATACCAGAGAAAATTCCATTCCCGTCGACAA tpg|BK006942.2|:138649-139981 7X4=65S 65S5=7X 
 tpg|BK006942.2| 251029 + tpg|BK006942.2| 251529 - INS GCCAATGGCAGTGGCGGCAATGTCAACAACAGCATCTCGTCAAATTCTACTTCTGACGACGAGATCTCTCCGTCGATCTACCAGCGCTCCAATTCGGACTTCCTGCCTAGTTCTAATTATGCTGCAGATTTCCAGTTTTCAAACAAGTTCCAGCCTCTCATGAGTCACCAGAGTCATAACGGAACCATTTTTCCAACCGTGGGCACCCAAAATGA tpg|BK006942.2|:250585-251973 7X7=100S 103S5=7X 
 tpg|BK006942.2| 62091 + tpg|BK006942.2| 62617 - INS CTGGATCAGAAGATGTACCGCTCTCAATTGGCCGTTTAGATGTACTTCCAATTTCTGTTATTTTTGCTCCATCGGTGCTATTGTTAGTTAGATCGGTTACGTTGGAAAAGTTAATCGCCGCTTTGACTGCAACTTCAGGTTGAATATTGAGTGTACGTAGGGGGGCATTCGTATTGATATTAGATTGGGATGCTGTGAATGGGTTCTGAAAACTTTGAAG tpg|BK006942.2|:61637-63071 7X5=105S 103S7=7X 
 tpg|BK006942.2| 312381 + tpg|BK006942.2| 312298 - INS TCTTGACGGACAAGCTTCGCAACTCGTTCGCAATGACCAAGTTTGGCTTTCGGGAAGCAAAGGGGAAAAAAATGAAAAATAAACTAATTGAAGTGGTAAAAAATAAGCTGTGTGTGTGCATATACATCGTAAGTGCGTTGGCTGTTCTGTGGAAAAGGGAGACACTTTTTATATCAGGTGCAAAGGCTTCGTACCAGCGTTGAAAAACTAAAACAATATTGAAAAATGAGTGAAGAAGGTCCTCAAGTTAAAAT tpg|BK006942.2|:311776-312903 7X62=1X161=14S 5S1=330S 
 tpg|BK006942.2| 242299 + tpg|BK006942.2| 242356 - INS GAACAAAAGAACTGTATGCCACCGGTGTTGACAATTTCATCAGTTTCCAGCAAGCAGACATCTTTAGTGGTGACTGGAAGCCGGGAAAGTATGACATTGTGTTGGATAAAGGGACCCTAGATGCCATTTCATTGAGTGGCATGAAGATCAACGGTAAACTTGATGTAGTCGATGTATACGCCGGAGTAGTGG tpg|BK006942.2|:241901-242754 189S91= 168=7X 
 tpg|BK006942.2| 135363 + tpg|BK006942.2| 135464 - INS ATCTACCTGCAGGAATCTAGACACTGACAAGTATTATCTCTGCTGGTCGGTACTTAAATTGGAGCTACAGAACAAGAAAGGTTAAATACAACAGATGGATTAAAGAACAAGAATTACAGCTGATGGAGAAATATAAAGGTGATAAAAACAAGGTAGCAGAACTTATTCACTCTAATTCTCATTATGCATTCAATTTAGTGGAGGCAAGGTTGCATCCAGCATTTGTGACACTTCTTCTCAGTAGCATTGGCTTTACTGCCTTTGGATGGTGTATTTCGGTGAAAACACCGCTTGCTGCTGTATTATGCACAAGTGCATTTGCAAGTTTATTTTCAAACTGTATTTTGACCTTCTCTACTACTTTGATAGTAGATCTCTTTCCGTCTAAGGCTTCTACCGCAACAGGTTGCTTAAATTTATTTAGATGTCTCCTATCCGCAATTTTCATTGCAGCACTGACCAAGATGGTCGAGAAGATGAGATATGGAGGTGTTTTTACGTTTTTGAGTGCTATAACTT tpg|BK006942.2|:134311-136516 7X307= 260=7X 
 tpg|BK006942.2| 429498 + tpg|BK006942.2| 429964 - INS GTGTTATTCTTCTTGTTAGCTTATTTGACAATATTCGCCATTGCGTTGGCCCTGGGGAAAAAGTGTGCACTTATAAGGTCGTTACTATCTTTATTGCAGTTAACAGTCTTCGTCATATGTATAATCATTACGCTGTAGGTTTCTTATTTTTATATGAAGCAGTGATATATAACATAATAAAGTTTCATCGCCTTTTACACAGTATATAGG tpg|BK006942.2|:429064-430398 7X170=19S 1S1=424S 
 tpg|BK006942.2| 300875 + tpg|BK006942.2| 301194 - INS TTGTTGATTGTCTTAGGAATGGAAATATTTAACAAATATACCTATAATGAAAAAAGGGTCCTTCTTTTTAATTATTATTGGCAGCGAAAAAGTTGTCCCAGCTTCTACTTTTTTTCCCGTTAAAAAAGGAAGCGGCGGAAGCTGATCTACTC tpg|BK006942.2|:300557-301512 7X76= 280S3=7X 
 tpg|BK006942.2| 32240 + tpg|BK006942.2| 32064 - INS TTTTTAGACAAGCCTTCATAACCACTGGATTCATAGACTTTTCTCCAACGCTCTGCTTTATGAAAATCGTCAAATGGGTTATGTGAAATACTCTCCGAATCTGATGTTAAGCTTTCTGCGGACACAGATAATTGGGCCTTTTCTACAATATCGTATTCTTCTTTTTGTACGGACATAGATGAAACTTTGTTTGTTGATTGAATTTTTTATTAATTGTTTGTACAATAAATAATTTCAATAATCAACAATTGAACGCTGCCTTTTTATACTAAATGATTCAGTAGAAGACGAACCTAGCGC tpg|BK006942.2|:31450-32854 7X265= 150=7X 
 tpg|BK006942.2| 325141 + tpg|BK006942.2| 325815 - INS TTTATCAACCATGCAAGCGAGAGGACAGCTGTTGAATCATCTGCATTCAATTGGATTGAAAAACGACAACACCAAGTGAGATCCGAAAACTTAATGAACAGATTATCTGCCTACTTTTTGCCCTTTTTGAGTAGAAGTTCTCACAAAGAACGTGTATTGT tpg|BK006942.2|:324807-326149 7X9=71S 75S5=7X 
 tpg|BK006942.2| 217943 + tpg|BK006942.2| 218167 - INS GTAGTTAACATGCACCATGCACCCTTTTTTATTCGTCTCTCTTTCCTTTTCTTTTTCCTCATGCTCTTTTTTCTTTTCTTCCTCATTTGGACCCTTTTCCTTCTTTGTCTTCTTTGCCCTTGCTTTTGCTCTTGCTGTCGTGGAAAGAACAGCTGTTGCTACCTTCTCTACCTCCTTACCACTTGCTTCCTCATACATCCTCGGATAACTGAATGCATCTTCTTTAGCGTAACAATTCATTTGAAATTTGGGTATAGCTTGATCGCTACCACGAATACCAATGACAGTTGTTGGTGTAAAAGAAAGGGATAAAAAGTGAGCCAGTGGGAACCAGTACCAGAATTGTGAGAACATGACCAAACC tpg|BK006942.2|:217203-218907 7X5=201S 11S341=7X 
 tpg|BK006942.2| 252493 + tpg|BK006942.2| 252332 - INS TCAGTGCTAAAATCTTTTAGAACTGTCCATCTTAGCCTTCCAAATTTTTCCAATTGTCCTTTCTCTTTAATTTCAATAACTGTGAACTTCTCTTGGTTCATTAACTCATTGAAATCAGACTCTGATAATTTCTCCAAGAATTCTATAGGTATATAGGGTGGGAAATTTATGATCTTCAGCTGCCACATACCTCTATTCGTCATTTGTTTTCTAAAGCTTTTCTCGTTAAAGATATGCTTTAATCTTTTGTGATTTATTTGAGTTTGTGAAGGTGTAATTGTTCCACCATTCTTTGCTTGGAGGGCACGGTCATCACCATTCGTACTTGTAGTG tpg|BK006942.2|:251652-253173 7X105=1X199= 167=7X 
 tpg|BK006942.2| 157390 + tpg|BK006942.2| 158037 - INS ACTATTATTCAGAGATAAAAGTACCGCTACTTGAACATAACAATAGTCAGCCATAATGGATTCATCAACGTTAACTTCGAATAAGTATGATTGATCTCTTGGCATGGTGGAAAATGCACATAAATCAGATGATCTATTGAAGAAGTGACCATAGAATCTACTCATTCTCAAACCTGTGGAACCACGGGCTCTCATTACGG tpg|BK006942.2|:156976-158451 7X152=23S 1S1=191S 
 tpg|BK006942.2| 318478 + tpg|BK006942.2| 319205 - INS ATCGTCATCTTCATTATCGTCCCAGGCTTTTTTTGAGTTAAACAATGGATCTGTTAACATCTTTTCAATTATATCGATTATACCGTTTCTCAGCATAAATGACTGTAAATTAGAGAACTCCACCACGAAGTTACAAATACTACCCAGAGTAATGCCCATAATCATAATTTCCGGTTTCATAAAATCTTGTCCAGCAAAATAGCATTCCTTGGTCAACGTATATGTTTTACTTAGTATCTGTAAAAGCAGCTGTGCAATTTTATTTCTCTTCAACGTCGTCCTAAGCGCTGAAACACTTCTCGAGAATGATTTCAACAATAGTAACCAAGCTGCCACGAAATCGTGATCATATATTGGGGGTAAACACATAGAATGACTTTCCGTAGTTGTTTCCTTTATCTCATCTTTCAAAGATATAAAATCCTGTAT tpg|BK006942.2|:317606-320077 7X175= 215=7X 
 tpg|BK006942.2| 147214 + tpg|BK006942.2| 147128 - INS GATGGGCAATACTTGATTCATTATTTTTCTTTTTTTCTTCCTGCTCCTGTCCAGCAATAGGAATTTTTTCTGATGTAGGAGAGAGAGATTTCTCATGTTCTAAAGATTCCAGATTTATGCTATAATGGCCGCTTTTGATTGCTGCCACATGAAACAACCCGACTATCTGTAAGCTACCTTCGTTATTCAATATGTAAACGAGCGGCAATCGCTCTATCGTATCAACACCGGAACAAGGTTCTAGAATAGTGCCTGAAGTAACGACGTCAACTGCCACACCTATTGGATTTGTGTCCTTATC tpg|BK006942.2|:146512-147830 7X222= 283=7X 
 tpg|BK006942.2| 178566 + tpg|BK006942.2| 178878 - INS ATTGATCGTCCTCAAAACGGTCGTCTCCCTTTGTTGAAGAATTGCGTCAGACACGCCGGGACATCTCCAAGTTTTTAGTGGACCCTGCGAATGGGTTTATCAACGGCAAGTACAATTATATTGTTGGGACACCCATGATTGCCGACACATTGAGATCCGGACTGGACATATCCACTTTATTAGCTGCGAACACCGTCCACGATGCGCCATCTGCTTCCCATCTTCCGTTCGATATCAATGACCCTGCCGTCCTGAACACGTTGCACCATTTGATGTTGCACATGCGTTCGATATACCCCATCAACGATAGCTCCAAAAATGCAACGGGTATTGCCCTGGGCCGGTATCCTGAGGACGTATATGATGGATATGGCTTTGGCGAGGGAAATCCCTGGGTCCTGGCCACGTGTACCGCTTCAACAACGCTTTATCAGCTCATTTACAGACACATCTC tpg|BK006942.2|:177644-179800 7X215= 426=7X 
 tpg|BK006942.2| 104198 + tpg|BK006942.2| 104352 - INS GTTTATATTATACAATTTTTTACTCCGTTGCAGGTCTCTTATTTTACATCCATGAGGCGCAATTGCCTGATAAGGATAGTGCTAGAGAATATTATGATATTTTGAAAGACGCAGAAACTGGTAGAAGCGTTCTTATTCAACTCAAGGATTCTAGTATGGCCGCTAGCAGGACTTATAATTTATTGAACCAAATTTTTGAAAAACTAAACTCAAAAACTATCCAGCTTACTGC tpg|BK006942.2|:103720-104830 7X160= 116=7X 
 tpg|BK006942.2| 274796 + tpg|BK006942.2| 274620 - INS TAATGGTACCACAAGCTTTTGAGCATCAATAGCCATCTTCGATTGCTTAATTGATTGAGTCTCTTGTTGAAGAGCCAGTTGAATGCATACTTTCAACACTTTTTTTTCTCGTTCATTTTTTCGCCTTATATAATAAGAATATTTATACATATGTAGATAATTTAAAGAAGTAGAAAGAGCCCTTAATGGTACCGCTTTACGAGGAAATTTAGCACTGTTACTTTTTGGAGAGTAGTGCAGTCTTAGAAGGGCCTTTGAGCTTGATGTACACGTCCG tpg|BK006942.2|:274054-275362 7X294= 138=7X 
 tpg|BK006942.2| 401874 + tpg|BK006942.2| 401713 - INS ACGTTACCATTCAAGTATGCAGGACTGCTGCAAGAACCAGGCTTGTAGCAGCAATTGAATTTATAAGAGATCTAAAAAACGAACATATTAATGCTTTTTGGTATAACTGCTCAACTGGAAATCTGATGCTAATTGGAACATTTGCTGCCCTGCTGTATGTGACTTCAGCTACGAAGGAAGAGGCTATGATTTTCAGAGATTATGTTAGAAATTATACCTGGGTATTGAAGATAGGTTCCAAATACTTTGATAAACTATCGAATGCTTTGAATAATATGCATTTACTATTTGCACAAATTCCTGGTCTTCTGACCGATGAACCGGTGGTCGTGAGCCCTAACTCTAACAT tpg|BK006942.2|:401001-402586 7X48=1X136= 328=7X 
 tpg|BK006942.2| 159674 + tpg|BK006942.2| 159484 - INS ACTGCACAACGGTACGTTGTGCAGATGCATATCGTTCATGGAAGTGGTGGCCTGATCAATTTGCTGGTGTAACTGTTCTTGAGCAGGGGTTAGGAATTGTTGCTGCCCCATGGAAGGGACTGCACCCTGTGGCGGCATTCCCATCTGACCATAGCTCATTCCAGCTGCAGCAGGATCCTGCGGAGGCATGAATTGTGCTGGCTGTTGTAGAGGGGTGGCATTTTGTCCATACTGGAGCTGAGCTTGTGGGTAAACACGTTTCTTGTGATGAGACATTTTGCAGATGGTCTCAGACTTATATATTTATGTCTGTTTCAATG tpg|BK006942.2|:158830-160328 7X368= 300=7X 
 tpg|BK006942.2| 228481 + tpg|BK006942.2| 228929 - INS GTTCTGCCTAACTCAAGAAAACAAGTCGAGTCGTGGTTACAGGATATCACTAACTTAAGAAAAGTCTATTCTGAAGCTCTTTCTCCGTCGTCAACCCTACAGGAGCTTGATCTTAACTCAAGCTTGCCTACGCAAGATCCAATAATTTCTGGCCAAAAAAGGAGACGTTACGATCTTG tpg|BK006942.2|:228111-229299 7X3=196S 89=7X 
 tpg|BK006942.2| 257936 + tpg|BK006942.2| 258383 - INS GACACGTACACAGGAGCAAAGTGAATAACGTCCTTCAATGATAGAGACTTATCCAATAAGCAGCACTGGTCTTCTAAGATCACCGCCTGTGCACTTTTCTACGGGCTCTTTTAATTGTATAACATGGACAGTGATCATTGCATTTTGCATCCATAGGCATACTATGGCTTAAGGTATTACTATCTATCGCGCCTAATCTCTGGGAGTTTTGAGGCCGGTTTCGGAATCTCGGTATCTTGCGATGGGTCCAAAACGGTGTAAACAAAGCAGGGGATAGCAGCGCAGGCTTCAACATCTCAAACC tpg|BK006942.2|:257316-259003 7X166= 152=7X 
 tpg|BK006942.2| 39624 + tpg|BK006942.2| 39863 - INS CTTGGACTTGCAAGCCAGTAGCTTCCAGGACTTTTGGTATGGCGTATGCAGGGCCCACACCCATGATTTCAGGGGGAACCCCCACTGTTTGAAAATCGATGTAGCGACCTAGCACAGGCAGATTTAACTGGTTGGCTACGGACCTGCGGGCTAACAAGACACCTGCCACACCATCGGAGACC tpg|BK006942.2|:39246-40241 7X3=88S 87S4=7X 
 tpg|BK006942.2| 96662 + tpg|BK006942.2| 97258 - INS CCACTGCAGAAGTACAGATTATACGTTCGTCGGCGAATAGTGGACGTAGTGTTACGAACGAACTGTATCGCGGATTAAGCATAAATTTGTTTGGAAATGCCATTGCATGGGGAGTTTATTTCGGTTTATATGGTGTCACGAAAGAATTGATATACAAGTCAGTGGCAAAGCCAGGGGAAACACAGCTTAAAGGTGTTGGGAACGACCACAAAATGAATTCGCTTATTTATTTGTCTGCCGGTGCTTCCAGTGGGTTGATGACAGCTATCCTAACAAACCCTATCTGGGTTATAAAGACCAGGATAATGTCTACAAGTAAAGG tpg|BK006942.2|:96004-97916 7X170= 302=7X 
 tpg|BK006942.2| 31018 + tpg|BK006942.2| 31488 - INS CCAGCCAGCTAAGTTATGAATACCCCTCATCTCTATGATTCCGGAAGCTAAAAGAGAGCCTAAAATTTGGAAAAGAGGTATAGCACACCAAAAGAAACTTAGGCGGAATGTGAGCTCAGCTCCAGTATAATAATATGACAAGTATAGAATATTGTCCGGGATGAACCCGCCCTGTAC tpg|BK006942.2|:30650-31856 7X10=78S 83S6=7X 
 tpg|BK006942.2| 317290 + tpg|BK006942.2| 316865 - INS GTCATCTACTATACACTTATGAGAATAAGCCTTTCCTACTATTTTGTATCATGACAACAGGGTTCTGTCGCTTTGAATGCGGCCTTTTACTTTGCCATATTTTGATAATGAAAAAACTTTCGAGAAATATTTACTAACAGGATCGAGAATTTTTTTCCTCATTTAAACAGGTAGAGTTATTCGTAACCAAAGAAAGGGTGCTGGTTCTATCTTCACCTCTCACACCAGATTAAGACAAGGTGCTGCCAAGTTGAGAACTTTGGACTATGCTGAACGTCATGG tpg|BK006942.2|:316287-317868 7X279= 265=7X 
 tpg|BK006942.2| 171793 + tpg|BK006942.2| 172396 - INS CGTAATGAGTGGCTGTATTGATGCTGTATTGATGAAGAACACATGCTGTATGTTATTCCACCACAAATCAAGCCTCTATCGAGGGGTGAAGTATTGGGGTGTACTTCTGAAAGATTAGATAAAGAACAATACGATGCCATGGTATTCATCGGTGATGGTAGACTTCATTTGGAGTCTGCAATGATACATAATCCGGAAATTCCTGCATTCAAGTATGACC tpg|BK006942.2|:171339-172850 7X217= 3S21=1X110=1X57=7X 
 tpg|BK006942.2| 222863 + tpg|BK006942.2| 223295 - INS GTCAACGCCTTCAGGGCCCATGTTTCTTTTTAATACTGTTTCAAGTATCTCTATGAGAACTCCTTTAGGTAAATCTTCCATATTCGACGAGATATCAATAAGTAGCGCATCCACGCGGCTATCTTGATACAATTCCGTTTTCTTCAATATGTCCAGAATCCTAGTTTGATCAGGCATCATTAAGGCACTTTCCAGATGTATAGTCAACGCCTCCAGGAAACATTCATGTAATGTATTTCTATCTTCCAATGATGACCCATCCTTAAATTCCGAGCTTTTCTTCATAACATTTATGCTATTAACCAACTCTTCTGACTTC tpg|BK006942.2|:222211-223947 130S76= 300=7X 
 tpg|BK006942.2| 194175 + tpg|BK006942.2| 194373 - INS GATTTATGTCATAGAGGTATGGTATGGTACTCATAATGAAATTTCCCCCAAATTAGCTACTACCGCGACTGATGAAATTTTAAATTTGTTCAAAGACGTCTGGCAGAAACATCAAAGAAATCTGCCCACAGCTGACAATCTTTTGTGCTACTTTCATAATGTCATATTGAAAAATGCAGAGGTGTTATGGGGGTCCTTTAGTCCTAGAGGAAGAAAGAAAACCGGTGATTTTCATGATAAACTCATTAGCATTCTATCATTCGAAAAAGTATCCTTGATATCTAAACCATTTTGGAAATTTTTCAAGAATTTCACCTTTAGTGTTCCGCTATCCATTAATGAATTTTGTCAAGTTACAATTAAGATGGCAAGCGAATCAGTTTCCCCAGCTATAGTAATCAATTTATGCTTTAGAGTTCTGATGTTTTACTCGGCAACGAGGATTATTCCAGCATTACAAAGAAAAAATGACAAACAGTTGCGCAAGAGTCGCAGGATCATGAAGGGATTGTATTGGTACAGTCCTTGCA tpg|BK006942.2|:193101-195447 7X5=182S 11S165=1X329=7X 
 tpg|BK006942.2| 100110 + tpg|BK006942.2| 100759 - INS GTGTAAGATACATATGGGTTCGACGACGCTGAATTTCAACTCAGAGAGGAATTGTTCACGTTTGCGTTTGTTGTTACGTCCATGGATGTCGTAGTAGAAATTTGGCCAGTGAGTTGAGTTCTTTGTAATTGCGGGGCGCTTTCACCTAAAATCGAGCTCGTAGCTTGTAAAGACTTTTTCACCTTCTGTGCTTTTATCCCCCTCGGGTCAATTGATGAAGATTCAGGAGCAGGTATTTCTCCAAATTTGGACATGTGCAATTGCAGCTGTCTTGTCAC tpg|BK006942.2|:99540-101329 7X232= 139=7X 
 tpg|BK006942.2| 240577 + tpg|BK006942.2| 241023 - INS GGGTTACCTTAACCGTAGGCTTGTTACCTTCTCTTGTTTCTTAAGAAGAAACTAGCCACGGCCACAGCGCCGGCTAGTACGCCTCCAGCGACGACAACACCCTTGAGTGTTTCCTTCTGGATCTTATCCTCTACCATACTCTTCAAAGCGCCCACCTGCTTGTTATTACGCTCATGCTCAAATAAAGTGTCTACATATCTCTTCGCCATAG tpg|BK006942.2|:240141-241459 25S87= 70=43S 
 tpg|BK006942.2| 234630 + tpg|BK006942.2| 234605 - INS ATCTTCTAGGTCATAAATTTTAAAAAGTCGAATTGCTAAAGATATTTGCTCAGCTCTGGCCATTTCTACAATATCGTAAGTTAAGCCGTCCAGCAATTTATCAAATTTTGATATTATTCCGGATAATCTTGAAAACAATTTCATGACTGTACGTTGTGC tpg|BK006942.2|:234273-234962 8X78= 157S4=7X 
 tpg|BK006942.2| 71609 + tpg|BK006942.2| 72090 - INS AAAGGTGACATTTTCTCATTTCCAAGGTTTATAGCGCTTTTCATGCTACTATTTGCTGAAAAAGCTGCACCACTGCCATGGCCACTGCCTCCATGGC tpg|BK006942.2|:71401-72298 19S32= 49=7X 
 tpg|BK006942.2| 277878 + tpg|BK006942.2| 278351 - INS ATCCCAAGATGCTACAGCCATCTATACTTATCC tpg|BK006942.2|:277798-278431 7X13=3S 11S6=7X 
 tpg|BK006942.2| 388797 + tpg|BK006942.2| 389499 - INS TCCTAAGAGTATGTAAGGTATCGAAATAATATCTTAATTTAAGAATGAAAACATCGTAATGAAGAAACGAACATGTTGGAATTGTATCATTAGAATACAACTGGAAGAGCGAGTAGCAACCACATAAAGTTTCCAAGAACCTTGATATTAGCAGCACCTTGGTAAGTACTCGAGATAGAAGGAACAGAGTATGTAGCGACTGCAGAACCAGAAGCAGATTGTAGTGGACCAGTTAGAGATGGAGATGTGACAACGGGAGCCACGCTAGAAGCAGAAGCTGTTGTAGCTAGTTGGGATGTAGTCTTGATTGAAATAGGGTTGGTTGCTGTGGCCACAGTTTCGTAATTCTTGGCACCATTTGAAC tpg|BK006942.2|:388055-390241 7X5=159S 5S348=7X 
 tpg|BK006942.2| 145855 + tpg|BK006942.2| 146109 - INS AAGATGTTTGCTCCTTGGTTTGGTAATATTTGTTGCAAATGCTGAAAACGGCGATTCGGATTTTGCTTTGACATGATTTCCAAATACAGGATTTTTTAAACCAGCCATGTCAATATTGGCACTTTTTTTTATAGTTTCAGTTAGCTTGCCTATGGGGGATTTTTGCGCTTCCTCCTCGACAACTTCACCATCTTCATCCGAGGGAGTTTCCGGTAATCTAGTAGAAGATGTTTGCTCAACCGTAGAATCTGTCAAATCATTACCGCTTACGTTGGGACCATTGCTTTCGTGTTCTTCATTATCGTCATTGATTTCACTGGTAGAGCCCTTACTTAAAGATCCATTTTCAGTATCATCTTTTGTGAAGGAACTGAATGGTGATTTGTTTCCTAACTGTGAAGAGAAAGGTGAAGCCTGAGTACCGAATTTAAAAGTTGTATCGGAACCAACAGATTCCAGAGCCTTTGAAAATCCAGATCCAAAGGAAGAACTCCCAAAATCAAAGGCATTGGTCTTTGGTTTCGTAGAGGTGTTAGGTTTCGTACCAAAAGGTGTCGAAGAAGAGTCTACAT tpg|BK006942.2|:144697-147267 7X198= 555=7X 
 tpg|BK006942.2| 426987 + tpg|BK006942.2| 427662 - INS TGCTTATATAGGAGAAGCTTGGTATAACACATGTATGACAGTAACTGTAGTTCTTAACGTACAACGATTGATATCTCATAGATTGAATACGGGGAGAGAAACACAAGAGAGCCCCATTTTGGATGCCAAAGAAAAGGATAATGGCAGCCATAGAGCCTTTGTCGCCCCTATAC tpg|BK006942.2|:426627-428022 7X10=76S 83S4=7X 
 tpg|BK006942.2| 248377 + tpg|BK006942.2| 248951 - INS TTGTTTTGCCCTGAATTCTGCGCCCCTCGGAGAAGTTTCTTTTCTTTTTTATCTCTTTTTCATCTCTGACCTTCGTTTCCTTTCATATAGACTACGCAGCAGAATCATGGCAGGAGCTATTAGCTGAGTGGGCAGATTACGTTTGCGCACTGTGCATTGT tpg|BK006942.2|:248043-249285 7X7=73S 71S9=7X 
 tpg|BK006942.2| 298004 + tpg|BK006942.2| 297673 - INS GGGTTTAACGTAAAGATAATTGATGTTGGTTTATAAGCTTCAGGAACGGATAATAAGTTCGATTTGAGCATGAATGGGAAAAAAATTCTAGTATGGAAGCCAAAACCTAAGACAATAAAAATCGCATAAATAAACATGGATAAGCAAAGCCTTGATAATTGAATACTCATCGGATGAATTAAACTATCATGCAAGATCTTAATATTAGGATCTTCTGGAGATCTGATAAAGAATAGAACACCTGGTCTAATGATATTTTTCCTAATCATTCCGATATATTTGGCAAACCAATACATGTAGAGAGTACCAATCGTCCAGTATACGAA tpg|BK006942.2|:297007-298670 8X8=201S 306=7X 
 tpg|BK006942.2| 371405 + tpg|BK006942.2| 371191 - INS GTCCTACCCTCCATGCTGCAATCTTACATAATTATTATATTGACCCCAAAACGGGCAGGGAAGTTGGCAAAGATGAAGAGTCCTACCCTAAGATGGTTTGGCCTACAAACTACTTCAAACTGGCGTGTCAAACAATGTTTACGTTATTCTTTGGTGGGAAACAATATGCTCCTAAGTGCACAATTAATGGAGAAAACATACAGGATTACTTGCAAGGAAGGTTTAATGATGCAATCATGACAC tpg|BK006942.2|:370691-371905 7X4=263S 228=7X 
 tpg|BK006942.2| 238861 + tpg|BK006942.2| 239451 - INS AAAAGATCAGGGATCCATAGAGCAGGGAACAAATCTCTTGCACGAATTTCTTCCTTACCATGTGTTTTTCTGATATCGACAAAGTCGAAGATATCTGCATGCCATGGCTCCAAGAAAAGGGCGAAAGCACCAGGTCTCTTGTTACCACCCTGGTCCACATAACGGGCAGTATTATTGAAAACACGAATCATAGGAATCAACCCGTTTGAAGTACCGTTGGTAC tpg|BK006942.2|:238401-239911 7X111= 6S3=7X 
 tpg|BK006942.2| 131714 + tpg|BK006942.2| 132340 - INS TTCACTGGCTTTGACTAGGACCGAGAGTGTAAAGCCAGAACCGGAGATAACCGCTCCGCCTCACTCACGCTTTTCCCGTTCTTTCAAGACAGTTTTAATAGCTCAGTGCGCTTTCACTGGGTTTTTCTCCACAATAGCAGGTGCCATCTACTATCCAGTTCTGAGCGTTATAGAAAGAAAATTCGATATTGACGAGGAATTGGTGAATGTCACTG tpg|BK006942.2|:131270-132784 7X217= 108=7X 
 tpg|BK006942.2| 198557 + tpg|BK006942.2| 198347 - INS AAGCTGTGGGTAGTAAACATTCTTGCTCGTTATAAGAAGCTGCGTCTAGTGCATCACTGGGCTGGGCTGGATCTTCCACAGTCATGCTAATTGGTCTTAGGTTGGAAGCACGAGTGTATTCCGAAACTTGTGGGTCCTCTTCGGGATTTGCCCCACCATAAGTGATCTCAATCCAGATGATGACATTGTTAACTGCTATGCGCAGCGGATGAAAGAGAAGCGG tpg|BK006942.2|:197887-199017 7X4=152S 26=1X183=7X 
 tpg|BK006942.2| 27129 + tpg|BK006942.2| 27461 - INS GTCTTGAATTTTAGAATACTTTTCTTTGGTGTCTCTGTAGCTTTCGGTTGGGTAAAAGGGTATTACTTCTTACTTCCACTGAAGGCTAGAATAACACGCAGGACTGAAAGGTGAAATGGCCTGTCTTGTGCTCTCTTCATTTTATTTTTTATTAGCAGAACATCCTGCTGTGATGAAATTTTATGGTCAACTTC tpg|BK006942.2|:26727-27863 19S82=3S 92S5=7X 
 tpg|BK006942.2| 235651 + tpg|BK006942.2| 236285 - INS GAAATCCCACACTGAAAAGCTCATACACGCTAGCTGGGTCATGTGCATCCGTTAGTAATGGAGGGTCTAGAGATAATACAAGAGTCCAATAGCCCACTATCGTGTTTATCCAGTACCCGTAAATACTGTCATACAAATAAAATATTGGCAGTCCAAAAAGCATATTCAATGCGACCACAGCTGCTCGAGGATCATAACAGCCCGACAGGATACCGCCTTGTATATCTCTGAATGAATATGAACCGGGAAAAAATGAATTGAATGCTACTGAAAACCCAGTGTTATAC tpg|BK006942.2|:235063-236873 7X245=15S 6S1=336S 
 tpg|BK006942.2| 168158 + tpg|BK006942.2| 168475 - INS TGGATGCTAGGGATTCATGATACTGGTTCAAAATTGTTGGTAAGTCCTGTATCGAGCCATTACCCAATGGCAAAAAAAACTTTTGTACTGATTTATCCTCCTGCGAGCTTGGTTGGTATTGATTCTCGATCGAAAAGAATGGGAATTGTACAGCATGTGATAATCTTAGTTGCTGTCTAACAA tpg|BK006942.2|:167778-168855 7X55=36S 6S1=259S 
 tpg|BK006942.2| 108748 + tpg|BK006942.2| 109476 - INS TGGTCAAACGTGGAAGTTAATGAAGTACATGCGGCAATCAAATATAGCTTCCATTGGTTTACTATTGTTTCCGGTAAAACATTTTTGAGTTTGAAATCAACATCATTTGCTACCCGCAGAATTATTTCGTGTACTTGCACAAGTCTTATACAAACGATAGATCGACACAATGCCATCGCCATAGGACAAGTTTTGAAAACCAACGCCAGTAATTTAGGAAAAGCCCTTTGCCATAGTGCAGCATCTACTCCGTACTCTGATTCGGCCAGTTTGATAAGTAGACC tpg|BK006942.2|:108166-110058 7X204=44S 10S1=286S 
 tpg|BK006942.2| 131002 + tpg|BK006942.2| 130904 - INS GGTATGCACTGCCTATTCTCATAAAAGCAAAAGTGCACAAAAATAATAAGGTGTGAAGCAATAGTAGAAAAGACACTGGGAACCCAAGGTATCTTATTTTAACAGATAAGTAAAACTAAGATCAAATCGCGTACTGATATCA tpg|BK006942.2|:130606-131300 7X4=67S 67S4=7X 
 tpg|BK006942.2| 306982 + tpg|BK006942.2| 307047 - INS CCTTCAAGTGATAAATTAAAGAGTCATTCAGAATCTTGATAAATATACCGACTTGAACAACGGGTCCAACTTCTAACCCGTCGACTTCTTTGGGCAAGTCTTCATGCGTCTTGATGAATTCGTCAAATTTCTCTTTTATTACTCTTGCTAAGAATTTGGCCACCGTGGATAGAAATTTGGATCTTTTATTGAATGAGGATGTTTTAAATGGGTCGAACTCTTCATCGAACATTAAACTAGAAATGATA tpg|BK006942.2|:306472-307557 7X5=119S 119S5=7X 
 tpg|BK006942.2| 428518 + tpg|BK006942.2| 429224 - INS GGAAGCAAAGTGTTTTCTTAAAAAGAAGAAATTACCGTGTTCTTGTGTTACCCAAAAATACTCCAGGATCTCTTACCATACATAGAAAGCATTCGGAAAAATGTTGAAATCGGTTAGCCAAGAATATCGATAATATGTCGCAGTAGAAGTTAAAGACAGATAGGAGAAGCTTGGTATAACACATGTATG tpg|BK006942.2|:428126-429616 7X4=90S 90S5=7X 
 tpg|BK006942.2| 213682 + tpg|BK006942.2| 213758 - INS GGTCATTGTTTGGATTTGAATTTAAGATGGAATTGTCCACTAGACCAGAAAAGTACGTTGGAAAGATCGAAACCTGGGATGCCGCTGAATCAAAATTAGAATCTGCCTTAAAGAAATGGGGTGGTAACTGGGAGATCAATGCTGGTGATGGTGCTTTCTACGGTCCAAAGATTGACATTATGATTTCTGACGCTTTAAGA tpg|BK006942.2|:213268-214172 7X12=13S 169=13S 
 tpg|BK006942.2| 294492 + tpg|BK006942.2| 294950 - INS TTTCTCCTCCCATTGTACGACAGCGATTGTGGTGGTTGATATTGATGATGTGGCATTTAGTAGTCCAACTAGGGGTATTCCAAGAACCAGCGCGACAAGCAAGGGATCAAATGCACAACTTCTCTCTAATTATGGAGATGAAAATAACCAGTCTCAAGATTCTGTTTGGGATGAGGGCAGAGATAATCC tpg|BK006942.2|:294100-295342 7X13=81S 88S7=7X 
 tpg|BK006942.2| 215818 + tpg|BK006942.2| 216255 - INS ATATTGCTGTTCTACAGTATAAGAACGGATTGTGAAGAACTCGGTGGAGAACATAGAAACAGACAAAAAATCATGGATTACTTTAATATCAAGCAGAATTACTACACGGGGAACTTCGTGCAATGTTTGCAGGAAATAGAGAAGTTTAGCAAGGTCACAGATAACACCTTATTAT tpg|BK006942.2|:215454-216619 18S23=53S 84S4=7X 
 tpg|BK006942.2| 112306 + tpg|BK006942.2| 112749 - INS ACATAGAGCCCAGTAGTTCGGCAAAAGAATTCCAATTCGAAGACTTAATTAAACTAGTTGATATAGAAAGTGGATCAGTAGTTTTTAACTGAGTAAAAACAATCTCTTCTAGCTTATCAGATAAATCTTCTTCTTCATTGCTGGAAGCCTGCTTA tpg|BK006942.2|:111982-113073 7X3=325S 78=7X 
 tpg|BK006942.2| 417351 + tpg|BK006942.2| 417731 - INS ATGCTTTACTTGCCTAGCGATTCCATTTCAAGAGAAAAGTTTTATTTAAAAAAAAATATCGAGGATTTTTCAGAAGACTTCAAGAAAAATCTTCTGTACATCAATGCGTTTGTTCTATGTGCGGTCAGCAACAGAACGACAAATGTTTGTACCAAGTGTGT tpg|BK006942.2|:417015-418067 7X5=75S 78S3=7X 
 tpg|BK006942.2| 69021 + tpg|BK006942.2| 69413 - INS ATGCATATTATATGCTGCACAAAACTCAGTAAGAATAGTTTTCAATTTTGGTCTTTTGATTGGTTTCGATAAAAATCCGTTCATTCCTGATTCCAAACATTCTTTAATGTTGCTATCGTCAGCAAAAGCGGTTAGAGCGACAATAGGTGAGGTATAACCTAAATCGCGCCTTATCATCTTGGTAGAAAGTAAACCATCCACTTTAGGCATCTGGACATCCATGAAAATCATATTATAATTTTCGCCCTTAGATGTCAATTCTTTAACTTTTTCGAATGCTTCTTGGCCATCGCAAGCC tpg|BK006942.2|:68411-70023 16S140= 69=87S 
 tpg|BK006942.2| 206491 + tpg|BK006942.2| 207046 - INS TATAGAGAGATCATACGTAATGATCTCCCACCAAGACCTGCCGACATTAACAACATCCCCGTAAAACATGATATTGAAATTAAACCTGGCGCAAGACTACCTCGACTACAGCCATACCATGTTACAGAAAAGAATGAACAAGAAATCAACAAAATAGTTCAAAAACTGCTCGATAACAAGTTCATTGTTCCCTCAAAGTCGCCCTGCAGCTCCCCTGTAGTCC tpg|BK006942.2|:206031-207506 7X104=63S 2S1=161S 
 tpg|BK006942.2| 59228 + tpg|BK006942.2| 59424 - INS CTATAAAATGTAACCACGTCAAAAAGTGCGGTAAGGCAACCACTAATGGTGCATGAAGAAATTTTGTTAATACATGTATACTGCATTGTATTGACGTCATGTTGATATGATTCAAAGAATCCAGCCAAATATTGAGATTGGTTGGGATATCATTGAAACTTGAATTTAAAGCATCGATATTCTGGAAGTAGCTTTCTGAACTTATTTGAACATCGAATGGAT tpg|BK006942.2|:58770-59882 7X3=201S 111=7X 
 tpg|BK006942.2| 406909 + tpg|BK006942.2| 406237 - INS GAATATATTGTTGTAG tpg|BK006942.2|:406191-406955 7X4=4S 1S7=7X 
 tpg|BK006942.2| 25886 + tpg|BK006942.2| 25364 - INS GAAGAAGAAGATTGACTGACAGAGCTTGAGACATCAGAAGTAGAGGAAGCTGATTGACTGACAGAGCTTGAGACACCAGAAGTAGAGGAAGCTGATTGACTGACAGAGCTTGAGACATCAGAAGCAGAGGAAGCTGATTGACTGACAGAGCTTGAGACATCAGAAGCTGAGGAAGAAGATTGACTGACAGAGCTTGATACATCAGAAGCTGAAG tpg|BK006942.2|:24922-26328 45S14=1X31=83S 17=1X89=7X 
 tpg|BK006942.2| 412538 + tpg|BK006942.2| 413088 - INS AAAATCACTTAAGACAACACCATGTTTAACCCACTGGTACAATTGACAACGTGATACTTCCGCAGTAGCGGCATCTTCCATCAAATGATTAATTGGGACACAACCAGATCCCCTTAACCAAGCCTCCATATATTGTAGGCCAATATCCAAGTTTACTCTGATTCCCTCAGTAGTGACTTGAGCATCTTGAATCTTCGTATTCAATAAATCAGATGATGTAACATGTACATCCGGGACAAAATATATTTGATTTGCTGTACCCATGTTACTGAAAACTTCATTACAAATCGGTGCCAATGCTGGGTGTGCTACCCATGAC tpg|BK006942.2|:411886-413740 7X163= 160=7X 
 tpg|BK006942.2| 219947 + tpg|BK006942.2| 220232 - INS TCTCTCTCACCAAGATTGTAATAAACTTTGGATGCAATCAAAGCAGCCATTTCACGGTCTGAAAAGGTATCGTCATCATACAATGCCTCAATATCCGGCAGTTCATTCGAGATCTCAGACCATAATTGGTCCACAACATTATTTATAGATTCTAGGGCATATGTTT tpg|BK006942.2|:219601-220578 13S99=19S 36S6=7X 
 tpg|BK006942.2| 331521 + tpg|BK006942.2| 331136 - INS GCTCAAAAT tpg|BK006942.2|:331104-331553 7X4= 5=7X 
 tpg|BK006942.2| 317867 + tpg|BK006942.2| 318162 - INS CTCTAAATTAATTGTAGGAAATACTACGAGTTCTGTGCATTCATTTAACTTTCAAAAGCAGGTCCATGTGATATAGTAACGTTCTGGCCTTTTCCCTGACAGATAATGATTCGTCTGTAATATTTTTTCTAACCAGATCGTATAATCCTACCTCCACGAGTTTTCTACATCTTTCCACCGTGGCACGTGTTACTTGTACATTTGATGTACTACCTTTTGCAGCCGGGGTGCGAACGAACTCATCGCCTTCATCATCACCCTCATCATTATCGTCATCTTCATCATCATTCGCATTGCTACTGCTATCATCGCCATCTGGCTCATCGTAGT tpg|BK006942.2|:317193-318836 10S162= 165=7X 
 tpg|BK006935.2| 699 + tpg|BK006935.2| 0 - INS CACACACACCACACACCACACCCACACACACCACACCCACACACCACACCCACCACACCCACACCCACACACCACACCCACCACACCCACACCCACACCCACACACCCACACACACCCACACCACACCCACACCCACACCACACCCACACCCACACACCCCACACACCACACCCACACACCACACCCACACACCCACACACCACACCCACACCACACCCACACACCCACACACCACACCACACACCACACCACACCCACACACACACATCCTAACACTACCCTAACACAGCCCTAATCTAACCCTGGCCAACCTGTCTCTCAACTTACCCTCCATTACCCTGCCTCCACTCGTTACCCTGTCCCATTCAACCATACCACTCCGAACCACCATCCATCCCTCTACTTACTACCACTCACCCACCGTTACCCTCCAATTACCCATATCCAACCCACTGCCACTTACCCTACCATTACCCTACCATCCACCATGACCTACTCACCATACTGTTCTTCTACCCACCATATTGAAACGCTAACAAATGATCGTAAATAACACACACGTGCTTACCCTACCACTTTATACCACCACCACATGCCATACTCACCCTCACTTGTATACTGATTTTACGTACGCACACGGATGCTACAGTATATACCATCTCAAACTTACCCTACTCTCAGATTCCACTTCACTCCATGGCCCATCTCTCACTGAATCAGTACCAAATGCACTCACATCATTATGCACGGCACTTGCCTCAGCGGTCTATACCCTGTGC tpg|BK006935.2|:0-2273 123S13=301S 122S561=7X 
 tpg|BK006935.2| 100744 + tpg|BK006935.2| 100956 - INS AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAGGTTTATTACCCTACTGCATTTTGATAATCTGAACATAATGAGCTAATGAAAGCAATTCTCATTTAAAAACAAGTATTCTCTCTTATTGAAGTATGCATTATCTATCATTATAAATTCTTTTATTCTGTTCGAGTCCATGTTTTTAAAAAAAAAAAAACATGTATGTATGCTCCATCTATATATGCTCCATCTGTATATTTTATATGCAAAGTTTTTTACAAGAGGAATTTGGGAACTGGAGGAAAGTGGCACAATACCTCATGTGGATAGTTCATTAATCTCTTCTTGTGTTAATGTGCTAATATAAAC tpg|BK006935.2|:100048-101652 7X310= 171=7X 
 tpg|BK006935.2| 29379 + tpg|BK006935.2| 28690 - INS TCTATCCTTACACAGAAATAGCCATAGGAAAGTGAATTTTGTCAGCCGACTAAAATTAAGGTTAGCTTACAAAGCAGCAAAAAATTTGACATCGCACGGTATTCCCTGAAAAAGGAGCAGGCAGGTGCTGTATATTTTTTTCGGTTCCTGCCTCTTACATGGCGTCGGTGTATCTTAAATACTAAAGTGAGCTGACTACCCTTTTGAGTGCCCTATGTGACCTCTGATCTCGAAAGTAAACAAGAGATACCTAATTTCACAGCCACTTTTTGTTGCGGACACTGACGGGATGTGTTGTGAATATTTTAAACCTTAAAAGTATTTATTGGTTAGTTATACTTAATTCTTATACGTCCTTTAAAACCAGTGTGCAGTAAGTC tpg|BK006935.2|:27916-30153 7X4=288S 369=7X 
 tpg|BK006935.2| 230216 + tpg|BK006935.2| 229775 - INS GTAGGATGAGTGGTAGTGAGAGTTGGATAAGATATATTGGGCAGGGGATAGATGGTTGTTGGGGTGTGGTGATGGATAGTGAGTGGATAGTGAGTGGATGGATGGTGGAGTGGGGGAATGAGACAGGGCATGGGGTGGTGAGGTAAGTGCCGTGGATTGTGATGATGGAGAGGGAGGGTAGTTGACATGGAGTTAGAATTGGGTCAGTGTTAGTGTTAGTGTTAGTATTAGGGTGTGGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGTGTGGTGTGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGTGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGTGTGGGTGTGTGTGGGTGTGGTGTGGGTGTGGTGTGTGTGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGG tpg|BK006935.2|:228603-230217 7X296=2I31=105S 9S4=387S 
 tpg|BK006937.2| 168159 + tpg|BK006937.2| 168810 - INS GTTTTGGGTCATCATGCACTGCTGTGGGTACGGCCCATTCTGTGGAGGTGGTACTGAAGCAGGTTGAGGAGAGGCATGATGGGGGTTCTCTGGAACAGCTGATGAAGCAGGTGTTGTTGTCTGTTGAGAGTTAGCCTTAGTGGAAGCCTTATCATATTCTTGAATTTTGGAAGCTGAAACGTCTAACGGATCTTGATTTGTGTGGACTTCCTTAGAAGTAACCGAAGCACAGGCGCTACCATGAGAAATTTGTGGGTAATTAGATAATTGTTGGGATTCCATTGTTGATAAAGGCTATAATATTAGGTATACAGAATATACTAGAAGTTCTCCTCGAGGATTTAGGAATCCATAAAAGGGAATCTGCAATTCTA tpg|BK006937.2|:167397-169572 7X7=270S 74S113=7X 
 tpg|BK006935.2| 30567 + tpg|BK006935.2| 30961 - INS TCTCAGAGAAGTACGTTTCGTCGCACAAGCTAAAATCATTGACAGGGCATGAGTTACGTCAATCTCTGGTCAATCCATGTCCAAAAAAATTTCTTGATTTGTTCAAAGTTTTTGCATAGGCACATTAATTGGTTTAGCGAAGTATACATTCTGAAGAACATTTTTGGGTGTATTTTCCACATAGAAAATTCGATTTTTTTTTTTAAATGC tpg|BK006935.2|:30133-31395 7X4=1X5=95S 99S6=7X 
 tpg|BK006938.2| 462562 + tpg|BK006938.2| 462513 - INS TAGGTTATTACTGAGTAGTATTTATTTAAGTATTGTTTGTGCACTTGCCGATCTATGCGGTGTGAAATACCGCACAGATGCGTAAGGAGAAAATACCGCATCAGGCAGTATAGCGACCAGCATTCACATACGATTGACGCATGATATTACTTTCTGCGCACTTAACTTCGCATCTGGGCAGATGATGTCGAGGCGAAAAAAAATATAAATCACGCTAACATTTGATTAAAATAGAACAACTACAATATAAAAAAACTATACAAATGACAAGTTCTTGAAAACAAGAATCTTTTTATTGTCAGTACTCTTTACATATGCCGCGGCTCGAGCGGCCGCATTTATATTGAATTTTCAAAAATTCTTACTTTTTTTTTGGATGGACGCAAAGAAGTTTAATAATCATATTACATGGCATTACCACCATATACATATCCATATACATATCCATATCTAATCTTACTTATATGTTGTGGAAATGTAAAGAGCCCCATTATCTTAGCCTAAAAAAACCTTCTCTTTGGAACTTTCAGTAATACGCTTAACTGCTCATTGCTATATTGAAGTACGGATTAGAAGCCGCCGAGCGGGTGACAGCCCTCCGAAGGAAGACTCTCCTCCGTGCGTCCTCGTCTTCACCGGTCGCGTTCCTGAAACGCAGATGTGCCT tpg|BK006938.2|:461167-463908 7X49=284S 641S3=7X 
 tpg|BK006935.2| 58922 + tpg|BK006935.2| 59282 - INS CAAGCTCCTCTGGTTCCTCCGCTAGTGGTTCTGTTTCCATTTTGATTTTCTTGCTATTAGCCGTTGGGCCATCGTTTCCAACTTCTTCATTGTCGTTGCCGTCGTCATCATCGTCGGATTTCCTCTTTGATGATGACGAGGACGGTACAGAATTGATGTACGTATTCATTAAATCCGTGTACCTCGAAGCAACGATAGACAATCCGGTGATCAGTTTCGTGCTGTCCATTTGCAAGATGGCCTCTGTGGACAGCTTGATAAGTATGTCATTGGGTAGCTGGGTCACATCCTGGTTGGAGTTCGAACTGTTCATCAATGAGTACACAGA tpg|BK006935.2|:58252-59952 7X280= 164=7X 
 tpg|BK006935.2| 3367 + tpg|BK006935.2| 3138 - INS TAGCTTGAACCTAAGTAGGGATATGTTTTTTTAGTAATTTCTTTGTAAATACAGGGAGTTGTTTCGAAAGCTTATGAGAAAAATACATGAATGACAGGTAAAAATATTGGCTCGAAAAAGAGGACAAAAAGAGAAATCATAAATGAGTAAACCCACTTGCTGGACATTATCCAGTAAAGGCTTGGTAGTAACCATAATATTACCCAGGTACGAAACGCTAAGAACTTGAAAGAC tpg|BK006935.2|:2656-3849 12S20=4S 205=5X2S 
 tpg|BK006935.2| 108741 + tpg|BK006935.2| 108773 - INS TCTCTCATCCTGTAGAAACGAAAATATTAGTGAATCCACCGGCCGCTTCCTTCTCGTCGTCGTTGTCCAGTTGCTCTGGCACCTTCATGAAACTCATAGAGATGACGTGCCCGTTGGTTACGCCGAAAAGGAACTGCAGTAGCATGTAACACAAGTCAACGATTACGGAGCCATTGTGCTCTTCATCGCCGCTTGAAGAGGAGGTGATGGCTGTGAACATCAAGAACAGTGGTATTGCGGCCACCCGCAACAATGAGT tpg|BK006935.2|:108211-109303 7X4=240S 129=7X 
 tpg|BK006935.2| 17805 + tpg|BK006935.2| 17954 - INS ATTTCAGCTTTTTGAAAACCCCATTTGGAAGGAATTAGGAAATTATTTTGCTTACTACGACCACTAATTTACCGCCATTTCTGGGCCTTTTTATTGACTATTTTGACCATGTGCTCGACTAGAAGAACGGCATCATAATCTGCTGGTAGAGTTAGTCTATAATGATTGTTGAAAATAAAGGCATAAGAGATATTCCACCTAAAATTCAAGTTATTGACTTTATTATCAGGATCTTAGTATCCTTTTTTGGTAAGTCATATTCAATGAACTAGGTCTCGCAAACTTTTTGTTCGAAAAGCGGTAGTGCATAGTTATGCTAACTCTGGATATATGGCATAAACCGTACAACACTAGCCCATTTTTTTGGAAGTAGTGAGGGCAGCTAG tpg|BK006935.2|:17019-18740 7X280= 193=7X 
 tpg|BK006935.2| 54925 + tpg|BK006935.2| 55336 - INS TTTAATGATGTCTTCCTTCAATTTTTCCAAATTGTTTATCAAGACAGATTGCGATTCGATCTTTTCCTTCAGTTGGGAAATCAAATGATCTTGTTTTTCTATAACGGAACTAGAATTTTCTTCCAATTCTAAGGAATCTAGTAGATGAGACTGCTCATTTAGTTTGGAC tpg|BK006935.2|:54573-55688 7X6=78S 80S5=7X 
 tpg|BK006935.2| 172810 + tpg|BK006935.2| 173055 - INS GTTAACGTCCTGATTTGTTTCCAAATGAAAGCTGCTGTCTTTGCGTCGTCGATAAAGGGAATGATGGTATCAATATTCCGGATAAAAGCAAAAAAAGCATCGTTGTCAAGCAGATCATTTAAAAAAGTGCTGTTTATATGTACTGTAAGGTAACAAAGCTTGGTGAAGTACTTTAAAACAGATAAATCTTTGATTTGGGCCATGTCAACAAAAAAAGATGTTAGCCAGGTAAAGAAACCCTCCGGTAATTCAATTA tpg|BK006935.2|:172284-173581 7X8=158S 240=7X 
 tpg|BK006935.2| 181623 + tpg|BK006935.2| 181744 - INS AACTGAGTACAATTTTGACGTATGCTTTCTTTAACGTTCACGATCGGGCTGGGCCATTAAACTTACCTTAGATATTATTTGGAACAGCACCGCAAGTGCTGATGTCCCAGAAATGGGCGCCGGTTCAATTAGGTCGTGAAGTCAGACATATGGAGACTCTCGGACTGAAAGCACTAAGGGATGATAGCTGGCATGCCAATTCCATTTTAAATTTACACATCAAGTTACAGGGTTTGGGAAAATCACGTTCAAAGCCTGAAAATTTGAGGTTGTTCACGGAAATCATTTGGTTATGTCTGTCGGCCTGCTATTTAGAGACATTTTTTATTGCAACAACCTACTCTATGCACTTACACGGAATCGCAGAATAACGCGCGCACAACACAATTGGGAAACGATAGGATTTTGAATAGTGTATTGCTT tpg|BK006935.2|:180763-182604 7X206= 397=7X 
 tpg|BK006935.2| 103238 + tpg|BK006935.2| 103531 - INS TAGCGTCACTACTCTTGGTGTTCTCTGGTTTTTCGGGAATTTTCTCGTATGTACCTTCCAGTTTCATTAATGCCACGGTTATTGGATCGTCATTAATTGAATCATCGAGCATATTAGCAATTTCATTTAAATTTTTCTTATTCAAGGAGCCTGTAAAAGCCGACTCAGAGTTTGCTCTCCGTGTGTTCCGGGCACTAGATGTGTCATTAATGTCGATATCGTCCATTGTCAATACACTTCCTGATATGTTACTATTAGTTTCACTCTCGTTCTTCAGAAATTTACTTTTCAGCTCTTCAAC tpg|BK006935.2|:102622-104147 91S9=112S 151=7X 
 tpg|BK006935.2| 45308 + tpg|BK006935.2| 45286 - INS TTGCATTTTTAAAGAAAAAGATAATCATTAATGCCTTCACGGGAATACGTATAGAACATTATTAAAAGTATATGAATGGCATATATATATAGAACACCACCCTTGGAAAACATTTATACCCCTTAAACTAAAACAATTTGCTGCGCTATACCGTGTTTCAG tpg|BK006935.2|:44950-45644 7X4=76S 78S3=7X 
 tpg|BK006935.2| 171256 + tpg|BK006935.2| 170677 - INS AACTGACTGAATATCTTGCAGTAATTCAAAAGTGGAAGGCCTGGTTCTTAAGTTCACATCTATCATTGAATGTATTATGGCATTAAGCCCTCTAGAGTAATACTCAGGGACGGTGTCACATTTCCCGTTTTTAATCTTAGTTTGTAGCTCGAGATAATTTTTTGCCTGAAATGGGGGGTGCAACGAACACATCTCAAAAATAACACAACCTAGTGACCAG tpg|BK006935.2|:170223-171710 7X4=156S 110=7X 
 tpg|BK006935.2| 62232 + tpg|BK006935.2| 62362 - INS GGTGGGAAGGGGTGGTATCCCTGGTATGTTCGTCTTTTTCGAAATGTCTCCATTGAAAGTCATCAATAAGGAACAGCACGGGCAGACTTGGTCGGGCTTCATCTTGAATTGTATCACCAGCATTGGTGGTGTCCTAGCTGTGGGCACTGTCATGGACAAGCTATTCTACAAAGCACAGAGATCGATCTGGGGCAAGAAGAGCCAGTAGAGGAAGAGACTGTCATAGGGAAGAGCCCTTTCTACATACT tpg|BK006935.2|:61722-62872 7X5=279S 124=7X 
 tpg|BK006935.2| 84081 + tpg|BK006935.2| 83893 - INS GGATACGTCTGAATGTATGACTTGGTTCTTGCTGTACATTCTTGGATTTCTGCTTTCGTTGGCAAAGGAACCGATAGTTCGAAATTAGACTGTCTCTTTGGAATAAAATCATCGAGCTTAACGTTTTTAGCGATTTGGTCAGTCAATATTGCCGGCTCAACGCGATCTGAGCTCAAAGCCGTCGAAACTCGTCCTTGAGAATGTTTTGGAGGTGGTAGTCTGTTAC tpg|BK006935.2|:83427-84547 7X156= 212=7X 
 tpg|BK006935.2| 5333 + tpg|BK006935.2| 5183 - INS CCTCCAAATATTCTAGAGGTAGCTTGTTGTGGTCACTAATGAGAACTTAAATAGTTTTCAACTGCTGGTGATAAATCAATAATTTATGTTCTTAACCTAACATTTGATGACCTTTGATGCGTTGGTTATGTTGAAGACAAATTGCCTCTAATCAGTTCCATTAAGAAATCTTCTTAACTCCTCCAAATATTCTGCCCATACGATACCTATTTGTTTACTTTGTCATTTTGCCATAAGATTGGTATCCACTTCTTGTCTGTAAAATAATTAGAAAGTAGCACAATTTTTACAGTAATGTAGCACGCGTAACTC tpg|BK006935.2|:4545-5971 7X8=165S 293=7X 
 tpg|BK006935.2| 197821 + tpg|BK006935.2| 197729 - INS TTCATCTGTTCCATAAATCTCGGCTTTTTATATACAGAACATTAGACGACGGGAAGAGAAAAACGTCAGTATAACCCACTTTTGTTCGTAAAAAAAGGTTATTCACTTCTACTCCGTACTAATCAATGACTTTAATGGTGAAACCATGATGAGGAGAGTAACAC tpg|BK006935.2|:197387-198163 7X93=30S 6S1=295S 
 tpg|BK006935.2| 135530 + tpg|BK006935.2| 135660 - INS GGAGTATAGCATCAAGATCGGTCTTCTCTGTTCGTGTCTTTTTCCTAACGTATATTTGCTTTGTTTCTTCACTCAACAATAAAGTCAAAGTAAAATTAAATACTAATTATTCTTAAAAGGGAAGATGCGAAATTTAGCGAAAATCTATTGATTATACACACAAAGGAAGAAAGGTAGTGGAAAGCTAAATAAAGGAGGTCATGGAGCCAGAGAGCATAGGCGATGTGGGGAACCATGCCCAGGATGATAGTGCCAGTATAGTGTCCGGG tpg|BK006935.2|:134978-136212 7X4=152S 135=7X 
 tpg|BK006935.2| 16471 + tpg|BK006935.2| 15802 - INS CTCCAGCAACATGTCAATAATTTTACTGGTGAGTAGCATTTATGACCAAAAGCGTACTTAAATTAGCAGCAAAAAAATTTTTAATAACGAAACTATAAGGAAAATACGAGGTACTGATTATGAGAGTCCCCGTTTCTCATTTTTGAGACATGATCTGAACAAGGCTGAAAACAGCAATCTTTTTCGATAACTTTTGCAAAAATTTCAAACATTGTTGTTTGAATGCAGCCAATTTTTATAGGGTACAGAGCTTAATGCTTTACATGTGCTTTATTTTCGGTAC tpg|BK006935.2|:15222-17051 7X6=160S 266=7X 
 tpg|BK006935.2| 146253 + tpg|BK006935.2| 146932 - INS GGAGCTGGTCTGGACCCATTACTTTTTCTAGCTTGGGAAAATGTACAGCGCCACCAAGATATGATTAGTGTAGATCTCAAAACTCCCCTTGTCATATTCAAATGTCACCATGGCTTTCACCAGACTTGCCTCGAAAACTTGGCCCAGAAACCCGATGAATATTCTTGTTTAATTTGCCAGACGGAATCTAACCCAAAAATAGTATAACATTTCTAAATATTTAATACAACTTTGGTTACATAAAAGTAAAATTTATACACCTCATTTCATTATGTAGATTCATATATAGAATACCAATTATGATTGACCCAATAGCC tpg|BK006935.2|:145605-147580 7X256=21S 2S1=21S 
 tpg|BK006935.2| 144846 + tpg|BK006935.2| 145006 - INS GGGTTGCGACTACTTGGGTGCATTGGAGTTCATAGAATCACTTTTGCAACCTTACTGTCCACTGGCAAACTTGTTGAAGCTAGATAATAATACGGAAGAGAGGACTAAGCAACTTATGGAACCATTTTACAATCTGTCCTTGGCTGCCCTAAGGTTTCTTATAAAAAAAGATAATGCCGACTACAATAGGGTTTACCAATTATTAATGGTAGTTGTTCGTGTTTTGCAGCAATCTTCCAAAAAACTAGACTCAATTCC tpg|BK006935.2|:144316-145536 7X204= 129=7X 
 tpg|BK006935.2| 117848 + tpg|BK006935.2| 118569 - INS AAGATAGACGCGTGAACGCAAGTCCTGGATTCGGTTGTTGATTGATATCTTGTGGTGCTGCTTCAATTTCAGCTTGAGTTTCTACTAAATTTTCAGGGACCATTGGATGATCAAGGTTAAATAAAACGCTACCAATAGTATTTGTAGAAATGGCAAAGCCCGCTAAAATGGGCACGGACTCAATCAAACCGGCCAAGAAACCAAATGAGGCATATTGGCC tpg|BK006935.2|:117394-119023 7X12=110S 14S193=7X 
 tpg|BK006935.2| 81542 + tpg|BK006935.2| 81121 - INS GTCTTGCTGAAAATTTTGTATTGCGACAGAAACCCGTAGGTGGCGTAGCGGTACCTTTTTCTTGATAACCCATTGGGCCATACAGGCTTCACGAACAGCACATTCTCTACAGCGCCTTTAGGCGTAGATCCCACTAGCACTGAAGAGGCCATGCGGGGTGAGCCATTGTGGCTAATTTTCGAC tpg|BK006935.2|:80741-81922 7X176= 92=7X 
 tpg|BK006935.2| 97137 + tpg|BK006935.2| 97359 - INS CTCTAGCTTCGCCACAGCCTCATTATAAATGCTATTCCATTCTTCATATTCTCCTTCAGAGATATCTCTCATCGCCAAACACAACGTCCGCAAACCCTCAGATGCATAATCTTCTAAATGTCTCATTGTAGCTTCTACATATTGATTAGCTTCATCATCCAATCTTTCCAGAATGACAGTATCAGCACCTTTACAGAATAACTTTATCGAACCATCCGGAAATCTAAATATAGCGCTCATTCTC tpg|BK006935.2|:96635-97861 7X13=10S 229=7X 
 tpg|BK006935.2| 88642 + tpg|BK006935.2| 89125 - INS ACTTTGAATTTGACTTCATCACTTAATCTTGAAGGTTTGTTACCTTTTATAGCAGCCAAACTTTGAATATGTGACTGTATTAAAGAAGATTGCTTCTTTTTTCTCTCCTTCAAGGCATTCTTCTTGTTTAAAGTATTCATGATTTCAACTTGTAACGTCTTCAGCTTGGAAATCTTATCATTATAACCATTTACTATCGTTTCGTACTCTTGCCTTTGCTTAGATGGAATATTTGAC tpg|BK006935.2|:88154-89613 7X226= 119=7X 
 tpg|BK006935.2| 176363 + tpg|BK006935.2| 176238 - INS CCGTCTTTCTACGGATACAAAAATTTATATTTATATACATGCGCCTAACTATTCATACTATTAATTTCATATTATTAAGCTTTTTTTTTTTCATTTATCATTTTTTTTCGTAACCTCTCATACCTGTACAGGTTTCATTCGTAAAGCAGGGACTCTAGTTT tpg|BK006935.2|:175902-176699 7X4=63S 141=7X 
 tpg|BK006937.2| 3114 + tpg|BK006937.2| 3856 - INS TAATAAACCTGCTATCAGTTGGCATCGAGAGCAAAACACATTGCTTTGAGATACCACAAGCTAAGAAATGCAGTGGCAGCAGGCATAATTACCATAGAACATGTTATCACAAAGAAACAAGTTGCTGACATATTTACAAAAATCCTTCCAGCTGAATCATTTAAAACACATAGGGCTGTCATGATAAGGGAACCAGAAACTACAAAATAACCATACTCATGCGTATTCAGTTATGGGGGGATGTTAAATGTGGTAACCTAATAGCATGATATGAGTAATGCTTTAGTATTGTTTCAGAGTTGTTTCAGTAATGTTTTAGACAAAGAAAACATATAATAGTAAACCTGTAATCAGGTAGTACTTAAGAAACTATACTTTCTGTGTACAAAACACTAACTATGTAATTCTTACATTTACATAACATGTAGAAAGGTCCAATAAACTTACTATATTATGACATATAAGTTAGATCGTAATTCACTACGTCAACATATCCC tpg|BK006937.2|:2106-4864 7X393= 10S472=7X 
 tpg|BK006937.2| 64696 + tpg|BK006937.2| 65304 - INS CTAAATGCCTCTTGCTTTACCATCCTCTCAATGTTCTCTTCTTTTTCCTGCTTATTTCTTAGGTGACCAAAAAGTGAAAAATTTTCCAATTTAACTTACGTCGTTCGAAGTGATGACAATAAGGATATTCATTTATTAATCGCTATTTGATACCCACTCTTGCTACTACCTCTCTTTTAATCCAAAATTACAATTTTTACGTTACCATTCATTACATAGTGTATCTCTATTCATTCAAGACTGTATTTTGTTTGATATATATATGTATATATACATATTATTTTCGTTAGTGTTCGGTTTCCAAG tpg|BK006937.2|:64072-65928 7X152= 168S3=7X 
 tpg|BK006937.2| 83132 + tpg|BK006937.2| 82937 - INS TTAGTATGTAGAAATATAGATTCCATTTTGAGGATTCCTATATCCTCGAGGAGAACTTCTAGTATATTCTGTATACCTAATATTATAGCCTTTATCAACAATGGAATCCCAACAATTATCTAATTACCCACACATTTCTCATGGTAGCGCCTGTGCTTCGGTTACTTCTAAGGAAGTCCACACAAATCAAGATCCGTTAGACGTTTCAGCTTCCAAAACAGAAGAATGTGAGAAGGCTTCCACTAAGGCTAACTCTCAACAGACAACAACAC tpg|BK006937.2|:82379-83690 7X121=15S 161S4=7X 
 tpg|BK006937.2| 20545 + tpg|BK006937.2| 20831 - INS GTGTGGTATAATTTAATGCTATCCATATCATCATCTCCATATTCGTCACTGTCGCTGTCGAGGTCCAGTGTTATGCATTTCGAGGAGTCAATTTCCCGTTTCAAATTATTAGCATAGGAGCTCAATAGTGGAACCCTTTTCTCATTTATTCTTGTCTCATCAGTTAGATTTAATTCAACACTTTTGTTCTCATGCAGTTCATCGTCATTCTGTACTGGTTTTGGATGTGCATTTTCCAGCTTTATATCATCGTCCTCATTTGAGGACGAATCGTCAAAATCAGCAAGAAAAGACTCTTTAGAAAAAAATTTTTTGGTTGGTATTGGCTTTTGCGGTTTTTTGTATTCGACATTTCTAGCTTTTTCCCTTTTAGAATCTTCTGAAGCCAATTCGCTTTGTATTTCCCGAATTTTTAATGTGTGTGGTACTTCATCTTGAAGTGTTTGTGCGACTGTATCTATTTGGGTTTTCTGTTCCTGATGCGTAGCC tpg|BK006937.2|:19553-21823 7X4=158S 245=7X 
 tpg|BK006937.2| 204504 + tpg|BK006937.2| 204942 - INS AGAATCCTTATCTCTTCATCGTATCCATTCTAGTTTTTGGATCAACGGAATGATTATTATAGTAGCGCTACCGGTAATGCAGTGAGTAGCTAGATCTATATCCAACGAGATTTTTTCATGGGCAACTCTAAAATTTCTAAACTTCATCTCATGCAAAGTGCTAGATTCACTAACAATGGCTCTAGGAGTGGCGTTTTTGGAAAAGGACATCATGAAGTCCACCTATTTATCCTGTTGTCACCTCTTCACTGTCCAAAAC tpg|BK006937.2|:203972-205474 7X295= 10S7=1X225=7X 
 tpg|BK006937.2| 170997 + tpg|BK006937.2| 171069 - INS ATGCTACGCCTGCATGACAAATAATGTTTGCACACGAAAAAAAAACCGCTTGTCCAGCGTATGCTACGCCTCCAAGATACTGTGCAGAAAAGACGACTTTTGGATTTAGTGGGTCTGCACGTATTAGTACCGCAACAATAACCATTACCAATGATATGAAAACAGAAACATGCCAATGCCTAGCTCTTGGGATCTTACTCATATATACAGCAGAACAAAGCGTAGAAACTATACCTACGGCAAATATCCCCGAAGGATAATTATTTCTTTGCGCCAACGTATATTTTTGGTTTTGTAACCATAATGCAAATGTAGAATTAGATGCGAAACCCAAGTTCTCACCTCCCAGAACCCAAACAAGAGAGAACATCCACC tpg|BK006937.2|:170233-171833 7X155= 8=1X343=7X 
 tpg|BK006937.2| 250490 + tpg|BK006937.2| 251173 - INS CCCATAAACCTGAGTGAAGGGCCTTCATAAACTTTTCTACTTGACTTTGCATTCTCTGTAGGGCAATATCGGTTCTCTTATAGCGACCACCGAGTCTGTGTCCAGAATGTTCCAAATACGCCCTAGCAATCAAACCTTTGTTGGATTCGGACGTGATACCGCCTCTTTGGATAATCTTGTAGACCTGGAAGTAGAAATCCTCATTGTAAGGGTCCTCAGTGACAATTTGAGACAACTGATATCTGGTGATGAAGTCCTTATCACGAGGAGTCATTAAACCTGAGTATTTCAAGATTTTCTCCACTTTGGCATGACGAATCTGCAAACGTCTTTGCTCTTCAGGCGACAAATCTCTCTTCGATCTGCGTCCACTTTGCAGAGGCATTTTAGTTGCGCCAACCACAGGGC tpg|BK006937.2|:249660-252003 7X163= 13S377=7X 
 tpg|BK006937.2| 25283 + tpg|BK006937.2| 25340 - INS ACTTGGAGATGCGATTGTTGCTGTGCAAGAATTGGTTTGCGTCACCTGTAATCTCACCACTACTGTATACCCGCTCCTTATATTCAATGGCTAACACTACTAGTTTCCCTATTGCTCCCCAGGCCCCGCCTAATTGGTCGTTCACTCCCAGCGATATTAGTGGGAAAACCAACGAAATCATCAACAACAGCAACAATTTCTATGATTCTATGAGTAAGGTAGAGAGCCCTTCCGTGAGTAATTTTGTGGAGCCTTT tpg|BK006937.2|:24757-25866 7X3=312S 128=7X 
 tpg|BK006937.2| 159524 + tpg|BK006937.2| 159156 - INS CTTGTCCTATACCGCCAGATATTTTCCACGGAAATTTTGAAGCCAGCTTCTTTGGATTTTCTGGATCTACGGCTAAATCATAAGCTAAAAAAACAGGCAAAAATTCGTTGTATACAATCAAATGTAAAGCCATAATAAAATTCACCGATATAGGGTAAAATACTTTTGTATGAAAAACGTGATGAAATATACTACTTTCTTTACAACCGTCTGGAGCTGTATCTATATTGGCATGCACAGCGTCTGTTGGTTCATGCAGAGAATATGTCCTAATCAGGCCTACAGACTGTCTTCTTGTTAAAATAGGATCAATCGATTGTATGCTTTCAGTATCATCGTCATTGGTAGTATTCACTAGGGGACTATTTTCATCCTCTTCACTATCTTGTCCTCGAATGCTGTTCACATTCTCATTACGGTGGTGAATGTTTTCCGAATCATCCTGAATGCGCTTTTGCCAGGGTCTTCTTTTCGGCTGTATACCAAATATATTCTTCTTAATAAAATCACCGACCTCTAAACCGT tpg|BK006937.2|:158092-160588 7X206= 263=7X 
 tpg|BK006937.2| 259998 + tpg|BK006937.2| 260720 - INS GGGTATATACAAGTCGGATGATGGGGAAGACGAAGTGTTCAGGTTTTCCACATCTTTTGCCAATTCTGCTGCCGAAGTCATCGCTGTGGTAGTAATTGTGGTGGTAGTAGTGGTTGTCATTGTATTGTTATCCGTGGACGTGGTGGTGTTATTTTCAGTGATCGAATTTCGATGGTTATTGGCAGCAGAATCGTCAGATAGACGGGCCACCAGAGAACCATCTGAAACGCGATACACTTGAGTAGTTTTGTTGCAGCCTGTGGCTAAGTATTCACCATCGTTACTG tpg|BK006937.2|:259412-261306 7X2=2I191=19S 3S1=419S 
 tpg|BK006934.2| 343987 + tpg|BK006934.2| 343558 - INS TATTACCTGTTGATCTAAACCCTGAGTATCCGCCAACCTATTACCACCGTGGGCAGATGTATTTTATTCTACAAGATTATAAAAATGCCAAGGAAGATTTCCAAAAGGCCCAAAGCTTGAACCCTGAAAATGTTTATCCCTACATTCAATTAGCCTGTTTGTTGTACAAGCAAGGTAAATT tpg|BK006934.2|:343182-344363 7X4=254S 91=7X 
 tpg|BK006937.2| 27288 + tpg|BK006937.2| 27415 - INS TTGCGACATAACTTGTTTCAACTTTTCAAGTGCGACTTTTTGTTAAATATTATGACATAGAAGAAAGTAGAACAGCCATTATAAAACAAAAGAGAAGTGAGAATACTATTAAGATGGCATTCCAAGATCCAACTTACGACCAGAATAAAAGCAGACACATCAACAACAGTCACTTGCAAGGGCCAAACCAGGAAACAATAGAAATGAAATCTAAACACGTATCATTCAAACCCTCTAGAGACT tpg|BK006937.2|:26788-27915 7X100=21S 1=223S 
 tpg|BK006934.2| 295682 + tpg|BK006934.2| 295427 - INS TACCTACCTACACAGCCCAGTACCACCCTCCATAGGCGCCAAAACTGTAATACCACCAACGCCCAGTCCTGAGATGATTCTTCCAATGAAATATTGATACCATTTGTCAATGGAGGCGATTTGGATGATGATCCCAATTGAGTAAATGACGACAACAGTCATCAGACCAATCTTACGTCCATACATATCACCGAGCTTTGACAAAACTATACCTCCGATAGCGCAGCCGATGTTGAAAATAGAAACCATCAAACCGGTTCTGACATCGGAAAGATAGGTAGTCCCGTTTGCACGGGTGCTGCCAAATCGCCTAATGAAGTCTGTTTGCCTGACAAAACCAGATATAGTACCAGTATCCCACCCAAACAC tpg|BK006934.2|:294675-296434 7X267= 13S339=7X 
 tpg|BK006937.2| 127890 + tpg|BK006937.2| 128415 - INS ATATATCAAAAAAAAAAGTAATCAGATTTTATTTTATTTCGACATTACCCCTCAAATATATGACTGGTATGAATGATAATAATGCCGCTATTCCTCAGCAAACTCCAAGGAAACATGCGCTATCTTCTAAAGTTATGCAACTTTTTAGAAGCGGTTCAAGATCATCTAGGCAGGGAAAGGCCTCATCGAATATCCAGCCACCTTCTAATATAAACACAAACGTTCCATCGGCGTCTAAATCAGCCAAATTTGGTTTACATACCCCAACCACTGCTACTCCTAGGGTAGTTTCTAATCCTTCTAATACTGCAGGTGTGAGTAAACCGGGCATGTATATGCCCGAATATTACCAGTCGGCATCACCATCGCACTCTAGTTC tpg|BK006937.2|:127118-129187 7X345= 368=7X 
 tpg|BK006937.2| 83862 + tpg|BK006937.2| 83872 - INS GCCTTCAGACGGTGTTAGAAGAATTTAAAGAGTATCTGGGCCGGCTTGCCAAGATGCAAACCGAATAAGTATTTCAAAGTTGCATTTGCCTTAGCCGTCCTGACACCATTGGCTATTTGGATATTTTATATTGACTTTCGTGTACATTGATCACATCGACTGTTCTATTGGCAAATGAACCACGGGCATTGACTATTTTTCAGGTTACTACTATATATTATTGTTGGAATAAAAATCAACTATCATCTACTAACT tpg|BK006937.2|:83338-84396 7X162= 10S230=7X 
 tpg|BK006934.2| 57277 + tpg|BK006934.2| 56525 - INS TGTTCAGAGAGGATATAGACCAATTTTTGCCTTCGGAAGTACCTTCGTTGGGGTCAGATCACCAGAATGATGGTGAGGATTCAGACACTGACAGTGACAACTTTTTGCAAGACCCTGAAGACGATGTGGATGAAGAAAGCACTGGTAGAGGTACAGTCACTACCACTTCCACATCCACTGAGTCAAGAGGCCGTCCATCTTCTTGTATCTTCGTGGCAAGCTTAGCAGCAGCCCTATCCGATGACGAATTATGTCTGTCGGTGACTGAAAATTTCAAAAAATACGGTGATTTGGCTAGAGTTAAAGTTTTGCGTGATAACGCAAATAGACCTTATGCTTTTGTTCAATACAACAACGATCATGATGCTAAACATGCTCTGATCCGCGCTCAGGGTACTTTATTAAATGGCAGAAGGTTGCGTTGTGAACC tpg|BK006934.2|:55651-58151 7X6=182S 215=7X 
 tpg|BK006937.2| 98743 + tpg|BK006937.2| 98775 - INS AAGTACTTCTTTTTCCACAAAAGAATCACAAACTGCTAAATCTTCTCTTCGAGCAGTTGAATTCAAATCTGATGACTTGATCGGAAAACCACCTGATGTTGGAAATGGCGCACATCCTCAAGAAAATACCAGAATATCTTCAGTAGTAAGGGATACAAAATATGTCTCCTAC tpg|BK006937.2|:98385-99133 7X124=26S 4S1=228S 
 tpg|BK006937.2| 123486 + tpg|BK006937.2| 123346 - INS TTGTTGTTACTACTTCTTGTAATTAACTTACTGTCGCATTCCAAATGGACTGCGAAACAGACACGAAACAATTACGAAAGTGACGACAGAGTAAATATTGTCATTAAAGAGAATGATGACCTCCGGGTAAACTGTGAGAATAAGTCTAGACCATTCGTTAAACTTCATCTTTAATTGAGAAGCATAGTAAAAAATAATTAACAAGTTAACACAACTATCTTGACCCATGCTACCA tpg|BK006937.2|:122862-123970 7X122=54S 1=160S 
 tpg|BK006934.2| 288996 + tpg|BK006934.2| 288296 - INS CAATTAAACCAGTTCTAACCTTAGACAAATAATAAGTACCATCGTGGTGCTTCATACCAAATCTTCTGATAAAATCAGTTTGAGCAACAAAACCAGAAATGGTACCAGTATCCCAACCGAAAACAAAACCACCGAAAGCAACCATTAAACAACAGATGGAAACTGTAACGTAGGCGGAGGCGGGCTTCTTTGGAATTTCAACGTAGTTATTAGATTCTTCGTGATTCTCGTCGAAATCTTTCATGTCATCTCTTTCAGCTTTGTTGGATGGAGTAGACAAAGCGGAATTAGAATCGGATTCAACTGGCGACAAAGCATCAGCTGGAGTATTTTGGACTGCTGTATCCTCTTGATAGGCAGCTTCTTCAGACATTTTTGGCAGATTTTATTGTAAAAGTGTTTCAAAACCAAACCTTGATAAGAGGCTTTGAATATATCTTTTCTTTATGGTTTCTCCGCTTTTTGAGCGAATACTATGAACGAGTTTTG tpg|BK006934.2|:287304-289988 7X455=15S 363S4=7X 
 tpg|BK006934.2| 11344 + tpg|BK006934.2| 11094 - INS GAGTCCAACCATATTCAACCCGGCTAATACGCATAGATGTTCTATAACAGAAATATGTAATGGATACTAACCTTTTTCTGTGAGTAACTTACTCTTTGCGTTACACCTCCATCTGACTCATAAAACAGGAAGACTCAGATTTATTAACTTTAGCATTTACGCCGCAAATGGTAAATGCTCCGGCCCGATACCCTGAAATAGCAACATGTACGAAAGAAGGTATTCAACTGAAGCCTTTTAGACAGACAAGACTATTGGATTATCAAGGCACTATATTTTACCACTACAGTAAATACTTCTGATAAGAACGGCATGAATAATCAAGTAGGTTTTATAATACTGGTATACAT tpg|BK006934.2|:10380-12058 7X260=1X83= 5S9=1X13=1X33=1X266=7X 
 tpg|BK006934.2| 488686 + tpg|BK006934.2| 489345 - INS GTGGTTGGGCCAGGATTCTCCCCGGCCGTTGATGAAATTGACCCGAACGACTACTTTATTATGGACTTTTCTTTAAGACTATACAATGTCAAAGCCGAAGTCCCTCTGTTCACTTCTGGCTTAACGTATATCAAT tpg|BK006934.2|:488402-489629 7X5=62S 62S6=7X 
 tpg|BK006937.2| 173649 + tpg|BK006937.2| 173913 - INS TTTAAGGTGATTCCACTCACTGATAGTGAATTTGGTAATCACGCCTTTAGCGGATTCATGTGCCAGGCCGTCTGTAATAAATCTGGCGATTAATCTTTGACCTTCACCATTTCTTGTCAAAACAACTGGTTCTTTAAATCTCCACGTTATTCTCTTCTTTTCTTTACTGAAGGAGCCCTGAGGTTTTGATAAAGCGCTTGTTGCATTAGCAC tpg|BK006937.2|:173211-174351 7X5=78S 186=7X 
 tpg|BK006937.2| 314460 + tpg|BK006937.2| 314082 - INS GCGTATAAATAGTTTGCATATTCTGGTCCAGCAGGGCAAGGTCCTCTATTTGGGTGTATCTGATACACCTGCTTGGGTTGTTTCTGCGGCAAACTACTACGCTACATCTTATGGTAAAACTCCCTTTAGTATCTACCAAGGTAAATGGAACGTGTTGAACAGAGATTTTGAGCGTGATATTATTCCAATGGCTAGGCATTTCGGTATGGCCCTCGCCCCATGGGATGTCATGGGAGGTGGAAGATTTCAGAGTAAAAAAGCAATGGAGGAACGGAGGAAGAA tpg|BK006937.2|:313504-315038 7X221= 265=7X 
 tpg|BK006937.2| 186176 + tpg|BK006937.2| 186251 - INS TGCATAGAATTAAGAAACATGGGGTATCCGCCACCTACACGAAGGCTTGGAGATAAGAAAAGGTACCATTATTCCAATAATCCTAACCGAAGGCATCCTTCCGCTGTTTATTCCAAGAATAGCTTTCCAAAATCAAGCAATAATGGATTTGTATCTTCTCCTACTGCCGATAATTCAACAAATCCGTCTGTAACTCCCAGTACTGCATCTGTACCTCTTCCTACAGCGGCACCTGGAAGCACGTTTGGTATCGAAGCACCCAGGCCATCTCGATATGATCCGAGCTCAGTCAGTAGGCC tpg|BK006937.2|:185564-186863 7X175= 281=7X 
 tpg|BK006934.2| 517268 + tpg|BK006934.2| 517744 - INS CGTCTTGAAGCAACAGACTATGCTACAAGAGCTTGGCCAGGTGGTGTTGGCGACAAAAAATTGGGTGCTAACTATGCCCCATGCATCTTACCTCAACGACAAGCTGCCAAAAGAGGGTACCAACAAAATCTATGGTTGTTCGGCCCAGAAAAGAACATCACTGAGGTTGGTACTATGAACGTGTTCTTCGTTTTCCTCAACAAAGTCACTGGCAAGAAGGAATTGGTTACCGCTCCATTAGATGGTACCATTTTAGAAGGTGTTACCAGAGACTCTGTTTTAACATTGGCTCGTGACAAACT tpg|BK006934.2|:516650-518362 7X97=1X136=30S 3S1=495S 
 tpg|BK006934.2| 374649 + tpg|BK006934.2| 374449 - INS GGTATGTCTTCGTCAATGACACAGTCGTTCTCCCAAAAGTCATGGGCGAGCTTGCTTAAAACGGCGGCAGCGTTTTGACGCTGCGCTCTACTTGAATCTTTCTCATTAATGTACTCGTTATACTCTTTAAAAGTTGATCCACTGAGAGATTGTGACTGCGATGTTCTACGTGGAGTATAGTAACTAGCAGGATTGAGCCTCCTGCACTCTTTGAGCCTCAATAGAGAAGCGATCTCCTCGGAGAGTTTTCTTCCCTTATGCTGGTGACCATCTTTAAGTTGTTTGTGTTGTCCTTGTGAAACTGCTGTTTCCATTTTGCCGCGTGGAGACATCTGTCCAAGTTGCCCCTGGCTCTCTGTAAATACCCATATATGAACGTTATATATATTGTATATTAATGG tpg|BK006934.2|:373633-375465 7X273= 140=1X60=7X 
 tpg|BK006937.2| 181400 + tpg|BK006937.2| 182050 - INS AATACCATATATTGGACCTGAACAACCATATATTAAGATTCGTCGAAGATCTGAAATCGCTGAGCGCTGTTCCGATTAATGAATCTGTATTTGATCCTAAAAAAAGTTATGTGATGGTTTCATTATTAGATCTCTCGATAGCTTTGAATGAATCGGAGGACATCTCAAAGTTCAAGAGCTCTTCAAAAGTGATTTCAGAGCTCATTAAAGGTAATATAATGTGTGCTCTTACGAAATATGCCGCTTATGATTTCGAAGTCTATATGAGCACATTTTTTTGTCACAGTACAGAATACAAACTGGTTTATCCAAAAACTGTAATGAACAATTCCAGTTACTTAGAGCTATCATTTATAGTGACACTC tpg|BK006937.2|:180656-182794 7X228= 354=7X 
 tpg|BK006937.2| 257774 + tpg|BK006937.2| 258425 - INS ATTATAACGTCATAGTTGAAATAGCGCACGAAAACGAACAGAAATGGCTCATTTATGACAAGAAAGATCATAAATATGTCTGCACATTTTCCATGGAGCCGTACCACTTCATCTCCAACTATAATACCAAGTACACAGATGACATGGCTACAGGCAGTAATGATACGACTGCGTTTAACGATTCC tpg|BK006937.2|:257390-258809 81S127= 162=7X 
 tpg|BK006934.2| 245245 + tpg|BK006934.2| 245964 - INS GACATACCTGAAGCTGCAGCTTCTCCGCCAAGCCTATTATCTTTTTTGAGAAAGAATGTAGGCAAAGATCTGAGCTCTATTGCCATGCCAGTAACCTCAAATGAGCCTATTTCTATTTTGCAGTTGATATCAGAAACATTTGAGTATGCTCCACTTTTAACGAAGGCTACCCAACGTCCTGA tpg|BK006934.2|:244867-246342 7X5=86S 87S4=7X 
 tpg|BK006934.2| 119031 + tpg|BK006934.2| 119545 - INS ATAGAAGGATGGTTCCATTAATGCATCTCTTGATTAATTTAAATTGCAAAAAGATTTACAAGTTTGCGAAAAGACTGCTTTATTTCCGCTTGGCCTGTGAGCTGTGTGTTCTCTCTTCTAATCCAGTAGGCATGTTGCATAAATAAACCTTATATTTGATGTTGTTTTAGAAATGTAATCTATATATAATTTCGTAGTATAAATATTTATAAATAAAGAAGTGAAACCATACCACTCATAAATAATGCGGGATGGTTGTCCAAGTTTGAAAGTAACTAAAGAACATAACTCGATGTCATATCAAACGTACTGGCAAATAAAATAAATCATTGGAGATGGATGAGTGTGGCGATAAGGCCCACGTGAATGTACAAC tpg|BK006934.2|:118267-120309 7X206=1X81= 14S350=7X 
 tpg|BK006937.2| 42520 + tpg|BK006937.2| 43050 - INS GAACTTTAGAGTGGAACATTAGGAATTATCAACAATGTAAATTTAATAAAAGTTAATTTGGAGAACTTAACAGACATTCAAGGTGGCTTGATGATCGCCGATAACGAATCCCTCGAGGATATTACTTTCCTGCCAAACTTGAAGCAGATTGGAGGTGCTATTTTCTTTGAAGGTTCGTTCAAAGATATCATGTTCGATAGCTTGAAACTGGTGAAAGGT tpg|BK006937.2|:42068-43502 7X4=108S 206=7X 
 tpg|BK006937.2| 133844 + tpg|BK006937.2| 133956 - INS GGGTATCTTACCACTTCGCTCATTATCTTACTAATGTAGTATGCAAGTGGCGAGTAATAGTTATTGGATCTTTCTTTTATGAAAATGATCCTTTCCAGAGCGAACGAGCTGAGACCTGTGAATGTAACAAAACCGAAGTACGTTAGTATAAAGAAGAACAGCCCCATTC tpg|BK006937.2|:133492-134308 16S71=4S 81S4=7X 
 tpg|BK006937.2| 96538 + tpg|BK006937.2| 96864 - INS TAGATTACCCACAGAATCGGATGATGATCTTGTCAAGGCCATTTGCAACGAGTTATTACAACTACAAACAAATTTTACTTTCAATTTGGTAGAATTTTTGCAAAAATTCCTGATCGCCTTGAGAGTCAGAGTACTCAATGAAGAAATTAATGGGTTATCCACAACCAAATTAAATCGACTCTTCCCACCTACAATAGATGAAGTCACAAGAATCAATTGTATTTTTCTAGACTCGCTAAAGACAGCAATCC tpg|BK006937.2|:96022-97380 7X5=154S 126=7X 
 tpg|BK006937.2| 232434 + tpg|BK006937.2| 232394 - INS GGTGAGCAACAAGGGTGGAATTTCTAAATTAATGATAATGAAGAGTAATGGGAAATCTTCTTCATATAGGAAATTACTTGAAAATTTCAAAAACGATAAATTTAATAGGAAAGGATGGATGGTTATGTTTCGGAAGGATTTTGCTAGGCTTATCAG tpg|BK006937.2|:232068-232760 110S94= 78=7X 
 tpg|BK006937.2| 143421 + tpg|BK006937.2| 143864 - INS AATATGCTGTTGCTATCACGAAGAAGAAGGAAAAATTGTCAAAGGATGAAAAGAATTCGAAAAAAAATAAAATTCTTAAAGATCAATTACGTTACCTGATAGAATTTTTCAGGACAAAGTCTGAGAGCAAGTTTCCCACCGGAATCCTAGAATTGGAAAGTGTAAAAGAAAATTACGGCGACTCCCTGATC tpg|BK006937.2|:143025-144260 7X4=180S 6S174=7X 
 tpg|BK006937.2| 113077 + tpg|BK006937.2| 113007 - INS GTCCATATAGCTACCAATTTAGTAGCTGTAAGATTAAAAAACTTATCCCACGAATTTGATGTAATAGAGAATTATCTGCGCTATATAGCTAGCACCAGTGAACATCTATTTACTGCTATTA tpg|BK006937.2|:112751-113333 7X179= 106=7X 
 tpg|BK006937.2| 184240 + tpg|BK006937.2| 184754 - INS AATAGGCAAGCTATAGAGCAAATGGTGACCCAAAGGTTTTCATTCAAAAGAATAGAGAAGCTTTAGAAAGTCCTTATGTATCAGCACATTTACATGAATGGATTGATTTGATATTTGGTTACAAACAAAAGGGGGACATTGCTGTGAAATCTGTTAACGTATTCAACAGATTGAGTTACCCAGGCGCTGTAAATCTAGATAACATTGACGATGAAAATGAGCGCAGAGCTATCACAGGCATTATTCACAACTTTGGTCAAACGCCTTTACAAATATTTCAGGAACCTCATCCGGAAAAAATAGCCTGCAATGTTCAACAGCTAACAACAGAGGTATGGCGTAAGGTTCCAATGAAGCCAATATTTGAGAAGACAATCTTTAATTTGAATGAAAAGAACAGGTCCGTCGATTATGTTATACACGATCCTAGTTACTTCGATTCATTATACTGGAGGGGCTTCGCTTTCCCAAACTTGTTTTTCAGAACGGAAGAATCGTTAGTGTCATTG tpg|BK006937.2|:183208-185786 7X221= 2S492=7X 
 tpg|BK006937.2| 131775 + tpg|BK006937.2| 131913 - INS AAATAAAAAACTACTCTTTTTTATTTCAATAGTTCTCGTTATTAGTAGGTCGTGCTCTTAAAAGATTACCCTTTCAGTAGATGGTAATGGGAATGGACGAGCCAGTACATATGAATTCTGCTTTGTAGCAACACCTGCATATGCGTTGTACCAAGCAATGAAAGCAACAAC tpg|BK006937.2|:131419-132269 7X54=31S 31S1=146S 
 tpg|BK006937.2| 115844 + tpg|BK006937.2| 116115 - INS CTTGAAGACCAGCATGTAGGAAGGTGATGATATGCTCCGTAAATAATTGGAAATATTGAGATATAATAACGATGACAATACTAACAAAAGTAATAGGTGAGCTCCGCCAATTGATTGTTTTGTTTTGAATATATATTG tpg|BK006937.2|:115554-116405 7X5=64S 63S6=7X 
 tpg|BK006934.2| 226667 + tpg|BK006934.2| 225992 - INS CTTTAAATGCTTTAAATGCGGCACCGGATGCAGCTAATTCGTTTGGATTGTTAGAAGCGTTCTTGTTCTGTGGACCAAGAATTTCGACTGATTCTGGTAAAGTGTATTCCAAGTTAGTGGTTAATTTTGGAGTAAATGATACACCACCAGTCAAAAGAACAGCATCGATGTCCAATGGGTCTAATTCAGCCTTGGCAATGACAGAATCAACGAAAGAGGAAAATTGGGCGAAGACCTTGTTAGCTACCAATTCGTACCTCATTCTGTTGATAGAAGCGTGATAGTCGAAACCATCAGCTAAGGAATCGATGGAAATAGTGGCAGAAGTTGCGTTGGACAAAGTCTTCTTGGTAATTGAAGAG tpg|BK006934.2|:225254-227405 279S12=46S 340=7X 
 tpg|BK006937.2| 230030 + tpg|BK006937.2| 229649 - INS GTTCCAACGCCAAGGGAAAGCTAACGCTATCCCAGATATATCATTGGATCCACGTTCACTTCCCTTATTACAAGCAGAAAGATGCTAGTTGGCAAAATTCAATAAGACATAACTTGTCTTTAAATGATGCGTTCATCAAGACTGAAAAGTCCTGCGATGGTAAGGGTCATTTCTGGGAGGTCAGACCGGGTGCCGAAACAAAATTTTTCAAAGGTGAAAATCGTGGTTATGAATTTGTAAAGGACTCCTTACAAGACATTGGGAAGTATTTTGAAATAGATTCTACAC tpg|BK006937.2|:229059-230620 7X4=202S 270=7X 
 tpg|BK006937.2| 77486 + tpg|BK006937.2| 77712 - INS AGATAACCACTGCCAAGCTGGAAGAAATGGCTAGAAGGCACTAAAAAAAGAGCCTCGCAGCGCAACTTAAGAACTGTGGACTACTAAGGAGCAGCAATCCGCTGGACGTGGGGGAGTTGAAAGTTGGCCGGATACTGCAACCTGCTTATCTATGACTCGATGAGAC tpg|BK006937.2|:77140-78058 7X5=78S 78S5=7X 
 tpg|BK006934.2| 430349 + tpg|BK006934.2| 430401 - INS CGTTTGAGTTAAGGCAGATATATTGACATTGTATTTTCTGCCGTACTCAGTCAAAATCAAATCTCTCATTTGAGATTCGATAGTGATCCATTGTTCATCAGTGAATGAAGGCCATAAATGGTACGATTTGATAGTGATCGTGGGGTCACTGAGTAGAATCATTTTGGCACTTTCCTCGTTCGTCTTTAAAGCTCTTAAAAGTAGTGTAAGTCTAGAAAATGCAGTGTACGATGAAATACGGTCTAACCAATCATCATAAATG tpg|BK006934.2|:429811-430939 7X222=15S 2S1=214S 
 tpg|BK006937.2| 213914 + tpg|BK006937.2| 214394 - INS TAATATATACCATTCAGAAGGGTTAGAGGA tpg|BK006937.2|:213840-214468 7X2=1X12= 10S5=7X 
 tpg|BK006937.2| 146135 + tpg|BK006937.2| 145867 - INS ATAAGGCATGACAAAGATAATATAAACGGAGAATGATAGGACATAAACCCATATGTTTTGAACTTGGCCTAATGCAGAAAAATACGAAGGAACTAACCAAAGCATAGCGATAGCGTACAATAAACCACCGAAAATATATTTAGGCCATTGTGTAATGCTTCTAGCTGAAAGTACAGCAGTGGATATGAGAAGCAACAAACATGGAACTAATGGCTTGCCCATAAACTTCACAGAACTCAAAGAAGCAAATAACATGACCGTACAAGATAAGGCGCCCCAAGGC tpg|BK006937.2|:145287-146715 7X199= 249=1X16=7X 
 tpg|BK006937.2| 125388 + tpg|BK006937.2| 125588 - INS CCTCATTTGCTGGTGCATCTATCTGCGTACTTGTGGCGTCCTTTACCGATGAATTTACATTCACACCTGGGGGTTTTTCTTTCACAAGAAATCTGAAGAATTTGTAGCATCTTTCACTACTATAAAAGTAATAGCGAGTACTCCATAAACCATTATCAAGTAAATATTGATTCATATTGTCTGTGATTGCTCTCCATTCTTTTCCCTTTACCG tpg|BK006937.2|:124948-126028 7X4=102S 104S3=7X 
 tpg|BK006937.2| 78566 + tpg|BK006937.2| 78321 - INS AAAAGGAAAACATAATAATTGCTTTGCAAAATGGAAAACAAATGACTTTGAAAATGGGAGAAAACAAAAATTATATAGGTAATGTTGAGTTCTTGATTTTTTTTTTGTTTCTGTCCTTGCCACAGCT tpg|BK006937.2|:78053-78834 7X3=1X8=3S 112=4X3S 
 tpg|BK006937.2| 5771 + tpg|BK006937.2| 5320 - INS ACACATTGGCTTCAATGGAGATGTGACTGCACGAGTGAGACATTATCTGTATTAGCTTCACAACCATACTCTGTTAGTAAGGAGCCATAGTCGACATCTGTCCAGCTCAATCGGGTATGATATTTGATATCCCCAAAATACATGGCTGTACCATGTAAAATGAGCGGTATATCGA tpg|BK006937.2|:4956-6135 7X4=201S 154=7X 
 tpg|BK006937.2| 246468 + tpg|BK006937.2| 246707 - INS CAGCAAGACAATATGACTACGACGGTACCCAAGATATTCGCGTTTCACGAGTTTTCAGACGTGGCAGAGGCCGTAGCTGACCATGTAGTCCACGCGCAAGACGGTGCATTGGCTCCAAAGAACGAGAGGAAACACTCTGTTCCCAACATCAGCATGAATGCACTGGATATGACGAGAGAGGCCTCTTGCAAAAGCACAGCATCTGCCGCGGAAGGGAAAAGTGGTAGCAG tpg|BK006937.2|:245994-247181 7X115= 250S3=7X 
 tpg|BK006934.2| 255940 + tpg|BK006934.2| 256287 - INS CCCTAACCATAGAGATTATTCTATGGCAGATTAAGGTTGCTGGAATGGACAAGGAAGTTACTTTCATAACGACTTGGGTGTGGCCTCTGACTGCAATCATGCTATCCTTCATACTAATTTTATTTCAGCCCTTTTTCATTATAATATCGTTACTGAATAAATTCTACAATGACAAGTTCGATATCGATAGGTTGATAATAGTGACATGCATAATCTTGTCCACACTTATTGCGCTGTTAAGTTACATAAATATTGGACCGTTCCAGTACACAAAAAATATTCTAACTAGATTGTCCATCGGAGGCGTCACAGTCATGGCTTCCCTATCTGGGTTAGCC tpg|BK006934.2|:255250-256977 10S166= 163=13S 
 tpg|BK006937.2| 203901 + tpg|BK006937.2| 204374 - INS GCTCAGGCGTATTTTTAACCAATCTCGGTACGCTGAATTCTAACTCCCATGTAGATTTTTCATCAAGCAAATCGACACATGGGACCCAATATGATGCAGAACTGCAAATCTCACCATTTGAAGTGTAAACGTTCCATAACCAGGGCTTGTCAGCATACACAGTATCGAATTTAATACCCGACTTTGGGTTTCTGATTTCATATTCAATTTGTAATGT tpg|BK006937.2|:203453-204822 16S99= 68=48S 
 tpg|BK006937.2| 8097 + tpg|BK006937.2| 8358 - INS ATCAAAAAAAAAAAAAAAAAAAATTGCTGTGACACCCCTTCAATGTGGTGTCTATACACC tpg|BK006937.2|:7963-8492 7X6=24S 26S4=7X 
 tpg|BK006937.2| 29207 + tpg|BK006937.2| 29475 - INS AAGTGCAGAACAAAAAGATACAGT tpg|BK006937.2|:29145-29537 7X12= 9S3=7X 
 tpg|BK006934.2| 248267 + tpg|BK006934.2| 247944 - INS TTCCAATGCAATTGGATCTTACCACGTGGATTTAAAGATGGACTCATTGGTATCCAGTGTGGTGTCCTTATTCGAAGTAGCCACTGGCAAAAAACCAATATACAAAATATTTGGGGGATCTCAAATCGAGAACTTGGCTTTACAAAACATCCAGGCGCGTCTAAGAATGGTTCTTTCTTATCTTTTTGCGCAACTGTTGCCGTGGGTTCGTGGTATCCCAAACTCGGGTGGATTGTTAGTACTTGGTAGCGCAAATGTTGATGAGTGCTTACGTGGGTATCTAACAAAATATGACTGCTCCTCCGCAGATATCAATATGCAAAAATGTAAAATCATCACACAAAACATAAACAATCAAAATCAGCCATTTCCGCACCTTTTCCTCTGTCCACTTTCAACCGTCC tpg|BK006934.2|:247122-249089 7X315=38S 195=7X 
 tpg|BK006934.2| 469410 + tpg|BK006934.2| 469285 - INS CAAGACTAAACCTGTTCTCTACGAGCTCTAGAATCATCAAACATGATGTTTCAACAAAAATGTGAAAAATTTACTGACTCACCTGTGTGTTCTCTACAAGAAGCACAACTGCCACAGGAAACTGCCAATGCGGATGTAAGAGGGTTTTTCCTCAGGGATAATGGCATACCCTTTCGCAGGTGGAATATCCTAGAAGCGAGTGATCCAGTCGACGCTTACAAAGAAATCTCCATAAAAAGCGAAAAGTTTTTCTGTGGTAGTGAAATAAATAATGAACTGGCTGCTCTTGATACGTTAGGGGCAATAAAGATTATACTGCGGCAGATTGAAAAGGAACCAAATGCTAATAAAGTCATACAAAGTTGGCACAGGGATATTGATTTTGTAAGGGTTTCTAATTTGAAAAGAGACTTATTGGGGGAATTCAAAGGATCGAAAACTACCGAAAATACAAACTCTATAAT tpg|BK006934.2|:468343-470352 7X176= 188=1X246=7X 
 tpg|BK006934.2| 129475 + tpg|BK006934.2| 130033 - INS GCTTATACATTTATTTATACGTTAATGGAGAAGTGAAGGTCGATAAAGTGGTTTATGAAAAGGAATAGGGTAGCCATTTTCATTTTTATGCATTTCTATGATGTCTAAACATTAGATGCATTCGTGAACTTTTTCTTGCAGACGAGATAGATGTAATTA tpg|BK006934.2|:129143-130365 7X8=71S 75S5=7X 
 tpg|BK006934.2| 289574 + tpg|BK006934.2| 289799 - INS GCCTTCATGATTCCCCAACATCGTTGAACCTGGCTTTTCGGTCCTAACTTTGCACCATCTAGGATGAGACTATCTTGACTGTTTTACTTTTACGCATCGCTAGAAAATACGTGCGCGTTGCCAAATCAAAATTCCCGCAAATTGATGCGGTAGCGTAGTTCTGTTCCAAAATGAAAGTGAAACAACATAATGTTCCTTCTAGTTTTCGTGTCTGAAAGCTAAACCTCAAAGTTGAAACTAAAGCATGATTCCCCACCTCCTTCCTAT tpg|BK006934.2|:289026-290347 7X172= 251=7X 
 tpg|BK006934.2| 285658 + tpg|BK006934.2| 285299 - INS GGACATGTATTCACCGGAGAATATATCAAAATTAATGTTCAAACGTGAATAAGTTTGGATATAGTGGTGGATGGATAACGAGCGAAACCTATTCCATATCTTAATGGCATTCTCATCCCCATTTTCTAAGTTTTTGAAAAAACTACGGGCCTCACCGCTAATCCCACACTTAGAGTTTCCGTTTATCTCTTCCTTGGCAAGGTCCATGTTGATTTTAACGTAGACGTCGAATAAATGCTGAATTGGCTGCTTTTGTAACGTCTTTTCATCGCCGTATCTCTTAAAAC tpg|BK006934.2|:284711-286246 7X333= 270=7X 
 tpg|BK006934.2| 193950 + tpg|BK006934.2| 194132 - INS GTTTTGCGCTCTTGTCATATGGGCAATATCTTTTTCTAGAGCAAGAACACCTTTATTGTCTGTATCATCCAATTTAGGGAAAAACCTTCTCAAAACCTCTTGTGTTCTTGCACCATGAGAATGCTTAAATAACTCGGAAGGATCAACACCGTATTCGTAACACAACTTGGTCCATGCTTTCTCTG tpg|BK006934.2|:193566-194516 7X10=82S 89S4=7X 
 tpg|BK006934.2| 227547 + tpg|BK006934.2| 227622 - INS ACCATGTAGGGTCTTCCCACACGATGAATGTAGGACTTGGAATCCACAGGAATATCGTAGTTTACAACTATGTCCACTGATGGAATATCCAACCCTCTCGCAGCGACATCTGTAGCCACGAGAATAGACCTCTTACCTGCCTTGAAAAGATCCAAAGATCCCATTCTCTGGTTTTGATTCAAATCACCATGTAGCGCAGTGGCACTAAACTCGAGCAAATTACATAATCC tpg|BK006934.2|:227073-228096 7X162= 216=7X 
 tpg|BK006934.2| 457879 + tpg|BK006934.2| 458326 - INS TACCGCTCCTCATCCAATTTCTTCTATAGAATATCCGTTTGCCTCCAGGAGTGAAGAAATGATAGCAGTAACACTGTGAAAGCGAGACTAAGAGAAACGACTTAAAGCTCGAAGACTTCTTGAGGATACGTTTATGTTTCTGTGGCTTCTTCTTCGCGGCGCGGTTCTCGCGTATAGGAATGTTCTAAGACAAGAAGGCATGAAGTTATGTTAACAGATTCTATATCTACTCGCTACGCATATATAAACGGATTCATCATTGAAACAATGGTACTTGTGGTAATGTGTACGACGATTTCAACCCGAATAAAAGC tpg|BK006934.2|:457237-458968 7X187= 157=7X 
 tpg|BK006934.2| 231465 + tpg|BK006934.2| 232080 - INS ATCGTCCACTTATCTAAAGACAGCTTATCAGCATGAAATCCAAAACGTGGATTTTCAGGGATGTCTTATCTAGTCACCGAACCAAAGCGTTTGATAGTTTACTTTGTAGGAGACTCCCTGTATCAAAGGCAACGAAGCATCTTCAACTGGGAGAACATTTCCTGTTCTTCCCA tpg|BK006934.2|:231105-232440 7X3=83S 82S5=7X 
 tpg|BK006934.2| 413293 + tpg|BK006934.2| 413808 - INS TATGCATGCCGAAGTTCCGCTTTCAGATCATTTATTTTGATGTTGAATTGATTTTCTCTTATGCTGTTGCTATTTTTTACATTATTGGAACTCTCCTCGGTGCTTCTGAGACCATTTTCGAAATTTTCACTGCAGACGCCATTTTTGAACTTCAATTCATCTAACTCGTCGATTAACTTTTTATTCAAACTCTTGTACTTCTCTAGCTCTCTTTGTGAAACCATTAGTGCCTTACTTGCACTGTCCATAGAACTGATACTTTC tpg|BK006934.2|:412753-414348 127S199= 247=7X 
 tpg|BK006934.2| 455969 + tpg|BK006934.2| 456417 - INS GAAGAAGAGAGTATAATAGGCTGGGTTCCACGCACGATCTACCGCTGCATAATGTACCTGAGTATAATATCTTCGAGAGGGCTCATAGGAAGTATTTTTATACTGGACTACTGAAAAAAACATTTTCTCTAAAATTCAATATGGATCCCACCGACAGCACTAAGCTGGAAACATTTCATCTTATTGCGTACTATACGGAAAAGGATATTCATCAAGGAAGTTTGAGGAGACCTTCAGAAAATCCTTTCTTCCATAAATTTCGACCTTCACAGAAACTATTAGAT tpg|BK006934.2|:455387-456999 12S163=45S 66S5=7X 
 tpg|BK006934.2| 322804 + tpg|BK006934.2| 322916 - INS ATTCTATACTTTATCCCCTCAGCATATACTGTAAATGCCGTGTTCATCAAGAAATGGGCGCATTACTACAAGAAGTTTTGATATTTTTTGTAACTGTAATTTCACTCATGCACAAGAAAAAAAAAACTGGATTAAAAGGGAGCCCAAGGAAAACTCCTCAGCATATATTTAGAAGTCTCCTCAGCATATAGTTG tpg|BK006934.2|:322402-323318 38S172= 1S169=7X 
 tpg|BK006934.2| 173696 + tpg|BK006934.2| 173406 - INS GTACAAGAAGCGTGGCAACAAGGTTATGACTCTCACGACCGTAAGCGGTTGCTTGACGAAGAACGGGACCTGCTAATAGACAACAAACTGCTCTCTCAACACGGCAACGGTGGGGGAGATATAGAAAGTCACGGACATGGCCAAGCAATTGGACCGGACGAGGAAGAAAGACCAGCTGAGATTGCAAATACGTGGGAGAGCGCGATCGAGAGTGGTCAGAAAATCAGCACAACTTTTAAGAGAGAAACGCAAGTGATCACGATGAATGCGTTGCCGCTAATCTTCACCTTTATCTTGCAAAATTCGTTGTCACTAGCATCTATTTTCTCCGTCTCACATTTAGGGACGAAAGAGCTAGGTGGTGTTACACTCGGTTCTATGACTGCTAACATCACGGGTCTTGCTGCTATTCAAGGTCTGTGTACATGTCTGGACACACTGTGTGCG tpg|BK006934.2|:172498-174604 7X189= 224=7X 
 tpg|BK006934.2| 417053 + tpg|BK006934.2| 417447 - INS TTCCCAATGGACGTGGTCCCACGGGTGCCGGGACTGTCCATTTATAGGAATTAATATTCAAAAGGTATATGTCATCGTCCATCAAACCTTCCTTATTGACTTTGTGTGTGTCACCGCCAAATACAACAAAGGCATTCCCGCATAATACAGCAGCGTGGCCTACCCTTGGTGGTGGTGTAGCTTCA tpg|BK006934.2|:416669-417831 7X4=88S 89S4=7X 
 tpg|BK006934.2| 238454 + tpg|BK006934.2| 238901 - INS GGCTTGTTATGGTGGCTGGGGTCTACATTCTGTTGACAAATCCACCGTGTTTGGTACAGTATTGAACTATGTAATCTTACGTTTATTGGGTCTACCCAAGGACCACCCGGTTTGCGCCAAGGCAAGAAGCACATTGTTAAGGTTAGGCGGTGCTATTG tpg|BK006934.2|:238124-239231 7X13=66S 74S5=7X 
 tpg|BK006934.2| 252686 + tpg|BK006934.2| 253454 - INS TGTAAAATTCTAAGCCTCGCTCAATGTTTTCCAGTACTTGGTCTATACATCTGATGACGAAATCGCGGCGGTAACTGTATAGACCGCCTAGAACTTTTGTTAATAAGGGAATATTTTGATAGCTAATCTTATGTGGTTTTGAAAACAGAGAAAACAGCACTTTCTGAATAGCTACATCGTCCCAGTGAGCTTTCCGAACCAACTTGACAATGTGTTTGAAGTCTAGGCTACTTAGTTCACTTCTAATTAATATGCGATAAAACTGTTGTTCAGGCGTTATTG tpg|BK006934.2|:252108-254032 7X188= 141=7X 
 tpg|BK006934.2| 304301 + tpg|BK006934.2| 304372 - INS CCTATATTATGAGGAAGTCATTGTTTTCAAGGATTTATTTCACGAATGTATTATTGGTTTGAAATTTTTTAAAGATCATAATGAAAAATTATCTCCAGAAACAACAAAAAAACATTTTGATATATCAATGCCCAGCCTACCGGTCTCAGCCACCAAAGATGCTCGTGAGTTAATGGACTATTTGGCATTTATGTTTATGCAGATGGATAATGCCACTTTTAATG tpg|BK006934.2|:303839-304834 14S193=10S 7S7=7X 
 tpg|BK006934.2| 436160 + tpg|BK006934.2| 436029 - INS CCTGAAGATTTATAGGATCCAGTGGCTCGATATTTTCTATGTGCTGTTCATATGACAGAGGTGGTTCGTCATCATCGAAAGGTGGAAATCTCATTCTTTTAAAATGTGTTCTATCTCGTTTTTCTCTCCTCATTGCTATCCAAGTAGCTGACCATTGGGCAGTATATACAGGCTCTATTACTC tpg|BK006934.2|:435649-436540 7X234= 92=7X 
 tpg|BK006934.2| 511749 + tpg|BK006934.2| 511987 - INS TCGCTCCTCTTGTAAAGTATGTATGTATTTTCGTTTTATTTAAACTCCAAAAAATGAATAATTGTTCCTGCAAATTTCTAGTTTATCACGTCTCATAATCACTGCTTATACCTCACCATTCCATTGTACTTTGACATATTTACCCCTCATCTATATATAATC tpg|BK006934.2|:511411-512325 7X5=178S 142=7X 
 tpg|BK006934.2| 508721 + tpg|BK006934.2| 509269 - INS TTTTATTCAAAAATTTACTCTTTTGGCAACTGTTTATAAGAAGAATAAGTCTGAGAATTATACTCGTATAAGCAAGAAATAAAGATACGAATATACAATATGATGAATTTTTTTACATCAAAATCGTCGAATCAGGATACTGGATTTAGCTCTCAACACCAACATCCAAATGGACAGAACAATGGAAACAATAATAGCAGCACCGCTGGCAACGACAACGGATACCCATGTAAACTGGTGTCCAGTGGGCCCTGCGCTTCATCAAATAATGGTGCCCTTTTTACGAATTTTACTTTACAAACTGCAACGCCGACCACCGCTATTAGTC tpg|BK006934.2|:508051-509939 7X284= 164=7X 
 tpg|BK006934.2| 462391 + tpg|BK006934.2| 462930 - INS TCTAGGTGTAACAATGGACCAAGATGAATGCAGAACAAGAAGAAAAGGCTAAGAAGGCTAACAACCCACAACACAGTATAACAAAGGATGAAATTAAGCAATACGTCAAAGAATACGTCCAAGCTGCCAAAAACTCCATTGCTGCTGGTGCCGATGGTGTTGAAATCCACAGCGCTAACGGTTACTTGTTGAACCAGTTCTTGGACCCACACTCCAATAACAGAACCGATGAGTATGGTGGATC tpg|BK006934.2|:461889-463432 7X156= 8S221=7X 
 tpg|BK006934.2| 182322 + tpg|BK006934.2| 183033 - INS CTATATTTTTGCCAGAAATCGACGCAGATGAGAAGTTGAAGTTTAGCGCAGGAAATTTCTACATAAATGATAAGTGTACTGGTGCCGTTGTTTCTCAGCAATGGTTTGGTGGCGCAAGAATGAGTGGTACCGACGATAAGGCTGGTGGTCCAAACATTTTAAGCAGATTTGTCAGTATTAGAAACACAAAGGAGAACTTCTACGAGTTGACTGATTTCAAATATCCATCGAATTATGAATAAAAAAATTTTTGTGGAATAGAACCGCGAATGCAGTCACTTCATCCATCAACTCATGTAAATG tpg|BK006934.2|:181702-183653 28S130= 40=119S 
 tpg|BK006934.2| 187044 + tpg|BK006934.2| 186456 - INS CCCTGTGGGGTGGAGATTATCTTGACCAAAACATACAGAGTGAAAATTGAGGCAACTAGCGTTGTAATGCCTATCAGTTTTTGGTTATCTTGAATAATTTGGGGTTGAGAACGCATTATTGCGTTTTGCTTCTCCAACCATAAGTTAAAGTAAGCTTGAACTGTGGAGTTCAAATGGTTAATCATGTCTGAATTCAGATAGACCTTGGACA tpg|BK006934.2|:186020-187480 7X5=290S 106=7X 
 tpg|BK006934.2| 76436 + tpg|BK006934.2| 76149 - INS TTTTGTGGTTCCATCCTTGAGGTGAAACATTTAGCAATATCAAAGTTGGTTTGGAGGTTAAAAAGTTATGCTTATTCAAAATTTTGACTTCATCCAGGTTCCAATGATCTTTGAAATGCCGGATTTTTTTACCGTTAAACAAATGTTCCTCTAATGCATCTAATAATTC tpg|BK006934.2|:75797-76788 7X204= 5S154=7X 
 tpg|BK006934.2| 223807 + tpg|BK006934.2| 224054 - INS GTATATGTTCAATGCTTCATCGCACCATTGACACAATCTAGAATAGCCGTAACTGGATTCATGCATGCATTAACCAAAAATTTAAATAATTGACCAAAGAGCATTTCTTGATAAGTGGAATGTTCTATTCCAAATTCCTTGGCAAATTTTGGTTCTGTTAATAATTTTACTAATGAGTTATTGGCTGCATCGTCCTCGACTACGGATTTTTTTTGAATCATTTCTTCCTCAGTCCAAGGCAATTTGGCAATTTTCATACCAGCCCACCCAGCATGATTGAAAACTCCTGCTTTATCCTGATAAACGCCATGAGAAATGACACCCTGAAATAAATGTGGTCTGTTTTTTGAATCTGTAAAGA tpg|BK006934.2|:223071-224790 18S285=1X61= 339=7X 
 tpg|BK006934.2| 453309 + tpg|BK006934.2| 453892 - INS GCATAATGCACTGGAAGGGGAAAAAAAAGGTGCACACGCGTGGCTTTTTCTTGAATTTGCAGTTTGAAAAATAACTACATGGATGATAAGAAAACATG tpg|BK006934.2|:453099-454102 7X3=46S 44S5=7X 
 tpg|BK006934.2| 497496 + tpg|BK006934.2| 497728 - INS GTAGAAGTCATGCAATTCTTGGAATCCAGCTTCCAGCCGGTCTTTGTCTTGAGACTGAGAATCTGGGTTCTTTAGGACGCTCTTTTTGGTGCCGTCCATCAATAACTTGAAGGAACCTGCTTTTATCGGAGTATTCTTGGACATTAGTCTGATTCCGCTGTCTAAGAGGTTATTAATCAGGATAGGGGCCTTAGCAGGATCGTTCAAAGCCGCACGCAAATTATCCTGATGTGAGTTTTCCGGTGATGGGGGTGCCGCAGTGTCGATGAACGCCTGAGACAGGAACTTTGAGTCCAGTACTTCAGAGACCAGATGTTTGTCTGCAGCGGCCACATATATGCCCAGACCATATGCTTTGAAAGTGATCGATGAGACACAACGTACACCCTTACCAATCAGCTCATATTGCGTGGAGAAGGGCCACTGTGGGGGGCCCATCTTCTTAGGGAACGCAGAGATGGATGCGTCCACTGCAACGCTGGTGGCATCCGCCTTTTTGATCTGGGAATCGTCATACC tpg|BK006934.2|:496446-498778 7X241= 63=1X195=7X 
 tpg|BK006934.2| 523725 + tpg|BK006934.2| 523841 - INS AGGTAAGTTGAAGGTCCTTCATACTGTGATCTGCAATAAACCACATGGCTACCGCACTTCTTGTCACTATCCTATGTGGAGAAAACCCAGAAAAAACTTTAAAGCGTGATTGAAATCAATAATTTGGCAAAGAACTAGAACCATACGCAAGAAAACCTTCCAACTTTGGCA tpg|BK006934.2|:523369-524197 7X4=221S 86=7X 
 tpg|BK006941.2| 589312 + tpg|BK006941.2| 589094 - INS TATATATATCTCCTCCTCTGGATCAAGCACTCTTTCTTTTCTTTGGCGGCCGTAAGATTTACCTTTGTCATTTTTCTTCTTCTTTTTTACCTTAAAGTTACTTGCTTCCCTAATCGCGTTCATGAAATCTTCCTCATCGTCTTCAGATATTTCACCGTAGTCCGAGAATTCTGCCAACAAAGAACTGTCTCGTTCGGAATTATATTCATCTTCGCTTAATTGTAGATCATGAGGTACATCCTCGTCATCATATTCCTCATCTTGAATCAAATGCTTATAGTCATCAATATTTCCGTATAGATGCTCTTCATCCTCATCGTTAACTTTACCCGTATCAGCGCTTTCTCGTTCAGCTGATTGATTTTGCTGTTCCTTTTTCAATTTTCCTGCTGCCATCACAGATACACTTGAGGGTTTCTTTCTCTAGCTTCAGATTCATTGTTGACTGGTGTTATTATACAC tpg|BK006941.2|:588156-590250 7X245=1S 434=7X 
 tpg|BK006934.2| 183904 + tpg|BK006934.2| 184613 - INS CAAATTATTGATAAGTTTGTTGCTTCCTCTAAAGTAAACTAGCTGGCTTCTTTAGCTAAAGAGAACAGTGACTTTATTCTTTGCCATGTGGAATTTGTATAAGCTCCTACGATGAAACTCTTTACAAAATTCCAAGCCTTAGCATTGTTACGAATAGGGTAGTCT tpg|BK006934.2|:183560-184957 7X121=23S 9S1=223S 
 tpg|BK006934.2| 324500 + tpg|BK006934.2| 324479 - INS AACCCATCCAACTACTTGACGAAGACTCCACGGAGCCTGAACTCGACATTGACTCACAACAAGAAAATGAGGGACCCATCAGTGCGTCAAACAGCAATGATAGCACTAGCCATAGTAATGATTGCGGTGCCACAATTACCAGAACAAGACCTAGACGAAGCAGTTCTATCAATGCAAACTTTAGTTTTCAAAAGGCTCATGTCAGCGATTGCACCATAGTCAATGG tpg|BK006934.2|:324013-324966 7X170=27S 2S1=230S 
 tpg|BK006934.2| 448939 + tpg|BK006934.2| 449631 - INS GTCATGACAAGAGACAATCCGAAAATCCAAACAACCTGATGAGGCAACTCCGGATGATACAGTTCGATACAGAAACACTTCCACAAGTCTTATCGCACTACCTCCAAATTTATCCAGAAGTACCTGAGAATAACTCAGCAAATGACGACAGCGACCCATTGATGCACGCGAATAATTTCAAGAATATGAATGCCATTCTTTTTGATGAATTAAGCAAAGAACGAACGGGAGCCTACCATGGATCCAATCTAGAACTATATACTCCAAAAAGCGCAATTTATCATTTAAAATTTGACATCAACATACCTTATCCATTGAATATTATTATT tpg|BK006934.2|:448267-450303 7X256= 41=1X277=7X 
 tpg|BK006934.2| 139490 + tpg|BK006934.2| 139831 - INS TATATCCTTGATCGATCTTTTGATACTGCTCCAAGGTTAATATATCAATACCGCTTAGACCAAGTCTTTCAGCAGTAGCGACACACTCACCAGATATGTGATGAGTCTCTCTGAATGGAACACCCTTTCTGACCAAGTAATCTGCCAAGTCGGTAGCTAGCATATCCATCGTGAGAGCAGCTTCCATCTTTTCCTTATTTACAGTTAAGGTAGAAATAACACCTGTGGCAATCAGCATGGAGTGCTCTACAG tpg|BK006934.2|:138972-140349 17S31=1X84= 91=42S 
 tpg|BK006934.2| 400487 + tpg|BK006934.2| 399846 - INS TCGTATCTCACCAAACTGAAGGTTGGTCACTATCCCATGACCAAACGCTGCCTTCATGAATTATATCTGCTAACTGCGTCACATTATTGACGTACGCTGAATTGCTTATTATTGGTGATAAACCACACGAAATATACTCTTTGATGTCCACGGAATTGAACAGCGAATCTAAGAATCTCCAATGGATAGATGATAAATCAGTCAGACCCTCTACAGTAGAGGGGCAATCTAATGTAGAGTTCCCCTGCTCATAATGAAAGACGTCATGAGGAAAAATATATGGAGCAGTAGTTTCATTAAAAAAATCGGTCAGCTCACCTATAACCAGTCTCTTCTTTTGTTCATATAGCACAGAGCCCAGAGTGGGCCAACCGTCAATGGACGATTTTCCGTAGATGTTCCAGGT tpg|BK006934.2|:399020-401313 7X6=105S 1S393=7X 
 tpg|BK006934.2| 495672 + tpg|BK006934.2| 496144 - INS CCGTTGGCCACATCGGGATGTTTAGAAATAGTTTTGACCAGGCCCTCCTTAAGATGCTTAAAATCTGTATTCCTTACGGGAGTTATCTTGGCTAGCATTCTCATTCCAGAATCCAGTAAGTCATCAATCATCATAACGGATTTTGAGTCATCACGTTTCAATAATCTAGCTAGATTCTCCTTAGGAGTCTTAGAATCATCCACATCAAGGAAATATTTATGTAAATAAGTTTCATTTAGAGTGTCTGAAACAAGGTTTTCGTCATTTTCAGCTAGATAAAGACCCAAGGCATAGACC tpg|BK006934.2|:495064-496752 10S158=61S 71S4=7X 
 tpg|BK006941.2| 179854 + tpg|BK006941.2| 180331 - INS CCTTTACAAACAGATTTTATAATAACGGAAGAGCTGCTGAAAAAAAAAGCAAGCTGCAACTGTTATATTTGCGTAGATAAACTTTACAACCGGTAATTGGAAGTCGTAAGTACTTAGTTTGACGTTTTCAGTACTCGTTAAACTACTCCTTAAATTGCTTTCTAACCTCTTCTTGTTTGTCTCTGTTGTTACTTGCTCTGCGGTGGCGAAAAGACGAGCAAAGGAGGTTGTATATATCACTCAACACGGAATGTATTACAGCTTTCTCAAATAAATGTAGTTGAAAAAGACCATTAATCGTGAGAATAGTTACTGATCAGGTGATGAGACGATAAAAACAGTAATTGAGAGGGTTTTCACGGGTAGTGGGCACAATGTTTGGATTAAATAAAGCATCTTCGACACCTGCAGGTGGGCTCTTTGGTCAGGCCAGCGGAGCTAGCACTGGAAACGCGAATACTGGGTTTTCGTTTGGTGGGACTCAAACTGGACAAAACACCGGCCCAAGTACAGGTGGACTATTTGGCGCTAAACCAGCCGGATCTACAGGAGGATTAGGTGCATCATTTGGTCAGCAGCAACAACA tpg|BK006941.2|:178668-181517 7X210= 293=7X 
 tpg|BK006941.2| 409150 + tpg|BK006941.2| 409147 - INS GTTGAGATACAGTTGGCATCTCAATATCGGAAGTGGAAGGTTCTGTCTCCTTCACTGTGTTCTCCTCTGTGGTGATTACGGAATTTATTGTTTCGTCGTCACTTTTATTTACAGTTTTTCCACCAGTCGTATCCGAAATTTCAGTAGTATCATCATCTTTAACAAGCTCATCAACATCCTGAGAACTGCTCTCATTCTCGGGTTCGTTAAAAGTCACGGATTTAGTTACACTTCCAGTTACATGTTGTGGAGTTTTGACACTTGCCCCTGATTTTCCATCAATCACAACTTCATTAGCTTCTCCCGTTGGTTTCGGCGCTTCCTTAATAGGTTCAGAT tpg|BK006941.2|:408457-409840 7X5=375S 169=7X 
 tpg|BK006934.2| 252188 + tpg|BK006934.2| 252806 - INS TAGTTTCTCTTCATACATTCTGCGTCAAGATCACCACCATACTCCAAATCAGAGTCGCTGTCTTCTTCTTCTTCATCATCATCATCCTCATCATCATCATCTTCATCATCATCCTCATCGCCTTCTTCTCCATCATCATCATCATCGTCATCGTCATCGTCATCATCCTCGTCATCGTCCTCATCGTCTTCATCTTCACTTTCGTCTTGCTTTGCCTGATGTTTTCCTGGCGCTGACTCTGTGTTCGGTGTACTTATCTCCGCGTCTTCATCTTCTCCTAGTAAATCGACACCATCGTCGTTTTCATCATCTTCATCCTCATCATCTTCGGTGATTGACTCGATAGGAACAGCACTCTCCTTACC tpg|BK006934.2|:251444-253550 7X135= 343=7X 
 tpg|BK006934.2| 387793 + tpg|BK006934.2| 387165 - INS AGTACCTTCAAGACAATCATCGACTTATTCTACCAACATTTAATAAGAACGTACCCAAGAATAAAAGTCCACAAGTATAACAATGTCTCGCGAAGGGTTCCAGATTCCAACAAATTTAGACGCCGCAGCTGCAGGTACTTCTCAAGCTAGAACGGCAACTTTGAAGTATATTTGTGCTGAATGTTCTAGTAAATTATCTTTATCCAGAACTGATGCAGTCCGTTGTAAGGACTGTGGTCATAGAATCCTGTTGAAGGCTAGGACTAAGAG tpg|BK006934.2|:386611-388347 8X8=146S 254=7X 
 tpg|BK006934.2| 390214 + tpg|BK006934.2| 390803 - INS TGTACTACTACTGAAGATGTTACTGGAACCTCTAGGGAAGAAACTCCATTGGCGGAGCCTACTAATGTTTCCAAAGAAGCTCCGGGCAATTTCCATATTCTGCCAATCGATCAAAGTGCAGACACAACCCAATCAAATGGTATAATTGGTGGACCAGGTCCTGTTCTTGTCCCAAACCC tpg|BK006934.2|:389842-391175 7X5=146S 39=1X50=7X 
 tpg|BK006934.2| 101475 + tpg|BK006934.2| 101220 - INS GGTTATAGGTCACTATCCTTTTTAGAGTCACCAGTCAAGGCTTTCATCCTTTTTTTGGCCTCATTTTTAGAGGCAGCACTTTCAGGCATGGCTGCAAAGCCAGGAACTGTATCACCTAAATCAATTTTACCCACGGAAGAGTTTCGTCTTCTTGTTTTTGCATTAACAACTAACCTATCGATAGATTTGTCCGTAGCTGATGTCATGTTGTCGTTATTTCTTCAGTTTCTCTGTATCTTGGAGTTCACTCTCAACACTGTCTAATATACCTTGCCACTTTAGATAGACAAGCAGTCAGATCAATTG tpg|BK006934.2|:100594-102101 7X209= 153=7X 
 tpg|BK006934.2| 282790 + tpg|BK006934.2| 282650 - INS TTAGGCACCACAATATTGGGTCCATTAAACGAAGTATTTTTCACTTGATAGTGAAAAATACTTCGTTTAATGGACCCAATATTTCGTCAACTTTACCGACTTGAGTCTTGTTTTCCAAATATATTGGCGCATTGAAATATGGAATCTTAGTGTTGATAGAACGGCAAACAATATCACCCTCACATGGATGTAGAAAAGCTCCCATTTCTAGAACAGTGTCTGGTGGTCCTTGTTGAAATGATCTAGCACTGCCTGTACG tpg|BK006934.2|:282118-283322 7X3=181S 17S218=7X 
 tpg|BK006934.2| 408242 + tpg|BK006934.2| 408974 - INS GGTTGATTATCTATTGAAGAGCACGTATGACCATCATTTTGAGAATACTAACGAAACGCCTATGGAATTAATGAGCAGGAAACTCCGTTTAGAAAGGGAAGCCTGGTGCTACTTTCAAGACAATTTTAAAGTCGGAAGCAAGACGCTATTCCACGT tpg|BK006934.2|:407916-409300 7X5=73S 74S4=7X 
 tpg|BK006934.2| 102183 + tpg|BK006934.2| 102191 - INS TCTTAGTCTAAGAAATTCGAATTACATAAATGAAACGCAATGGATTCTAACTGTTAAATATAGGGGCCATGCCAGAGGCAATGCGTAAATCTATCTAAGGAAACCGTTGACAAAAATGTCATCATCTGCGATTAAAATAAGGAATGCACTGTTGAAGGCAACAG tpg|BK006934.2|:101841-102533 15S29=45S 78S4=7X 
 tpg|BK006934.2| 235296 + tpg|BK006934.2| 235536 - INS TTAAGTTCATCCACTTCCAGCCTGGCCAAGTAGTCTGTGATGTTTTCGCCGGCGTGGGGCCCTTTGCTGTACCTGCGGGCAAGAAGGATGTCATCGTTTTGGCTAACGACTTGAATCCTGAGAGTTACAAATACTTGAAGGAGAACATCGCATTGAACAAAGT tpg|BK006934.2|:234956-235876 7X6=13S 143=7X 
 tpg|BK006934.2| 43448 + tpg|BK006934.2| 43679 - INS GTTGAGATCATGCAACAAAAATTCCCTGCTACAAATGTTACCACTATACTTGATGAGATCTTTTCAGGTTGCGACTCTACAAAACCCTCTCTGAGGAAGGCATCTTGTATTTGGCTGTTATCATATATTCAGTACTTAGGTCATTTGCCAGAAGTAAGTTCCAAATGTAATGATATTCACTTGAGATTTATGAGATTTTTGGCAGACAGAGATGAATTTATACAGGATTCCGCCGCTAGAGGGCTTTCTTTGGTTTACGAAATTGGTGGTT tpg|BK006934.2|:42892-44235 7X3=202S 136=7X 
 tpg|BK006934.2| 333775 + tpg|BK006934.2| 333905 - INS TCCCTAGGAATGAGAGGCAGACAAGAAAAGTGTCTATGCTGTGGTAAGAATCGAACGATAACAAAAGAAGCCATCGAAAAAGGTGAGATCAATTACGAACTGTTTTGTGGCGCACGAAACTATAATGTATGCGAGCCTGATGAGAGAATCAGTGTGGACGCATTTCAGCGTATCTACAAGGA tpg|BK006934.2|:333397-334283 253S53= 171=7X 
 tpg|BK006934.2| 166434 + tpg|BK006934.2| 166434 - INS ACCAACTTCTGATTCATCAATTTGCAAGAATGCCAGGTAATCACCAGTTGGTGACCACCACGCAGCCTTGTCGTCTTCAAAAACTTCTTCCTCGTAAACCCAATCTGGCTTACCGTTAAAAAGAAAGGAGCTTCCGTCGTTGGTCACAGCCCGTA tpg|BK006934.2|:166110-166758 7X23=1X113=8S 3S1=132S 
 tpg|BK006934.2| 474357 + tpg|BK006934.2| 475005 - INS TCTATGCTGGATTGAACTCAGGAAATGTTGTATTCTGTATCTTCCCGCAATCTGGTGGTATCTTATTAATTATCTCAGCAATCGGAGAGCTTCGAAAGTTGTTCATTTTATTTAGCTTCGATGTTTTAGTCTCCTTCAGTTCCGGTGCGGAAAGCTGTGTGTAACCTTGATTCATTTCGATAAAATTTGCGTTTTTATAAAATTCCCAAAAATACTGACTATGGTAGAAAAGATTTCAACGAGGAAGGTGGTAAAGATCAATGAAGTATCTTCAATCATTATGTAGGTTATAAGTAAATGTTTTTGTTTTCAAT tpg|BK006934.2|:473715-475647 7X9= 157=7X 
 tpg|BK006934.2| 125773 + tpg|BK006934.2| 125831 - INS GTGTATTGGAGAAAAAAAAAAAAAAAAAAAAAGGAACAATATAACTTTTGTAGTACGTGTGCCAGGTTACAGATATGGTTTCACTTCTATGTCGTGCTTTTTTCATTCATACGTAATCTTATGCATGTAGGGGATAGACGCACAAAAGCACCAAGGCTGCATGTATTGATAAATTGGCTTACACGATTCCAGCTAAGGGGACTCGGACGGAACCGTCTCATATTATACGTTCAGTGAATATTTTTCACGGAAGAATGG tpg|BK006934.2|:125243-126361 7X367=1X47= 242=7X 
 tpg|BK006941.2| 120597 + tpg|BK006941.2| 121268 - INS CTGTAAATCACTTGGGAGTTGTTATTGACTGAAATGCAAGATAAATAACGTAATGGGGTGATGTATGATATCGTATAAAACACAAGAAAGGATAACAGCACTATCATGCAAAATTGCTTATTTCTGGTATATTCTGGATTCCGAATGACACTTCCCTTACTGGAAAATCGAATTCAAGTGACCATTTAAATGGTCACCTATTTCTCAGGATGACCGCTAATTCTTCTCATCAGGGTTTCCCAAGTTGTTAGCAAACTGTATTGATATCTTTTTGCGGGAGTGAAACCAACTATTCAGCTCAGTATCGGATTAATCTCTCCACTTAATGCTACGGAGTTCTTCCAAACATTAGTACTGGTGCCAGTATCAGCACCACATCAACAGGTGAACTCAAAATTACATTAGTCAGGAGCAGTACACCCGTTAATCGTGGGAATCTCTGTAC tpg|BK006941.2|:119693-122172 7X244= 418=7X 
 tpg|BK006934.2| 514923 + tpg|BK006934.2| 514200 - INS GCCTCTCTACACTTCTGCCGCTCTCAAATTC tpg|BK006934.2|:514124-514999 14S98= 16=7X 
 tpg|BK006934.2| 286412 + tpg|BK006934.2| 286215 - INS AAATTCTACTAGGTACATCATGCAGTGCTTTTGAGATGTCTAGGCG tpg|BK006934.2|:286109-286518 7X11=17S 15S3=7X 
 tpg|BK006941.2| 298675 + tpg|BK006941.2| 299341 - INS GGTTTAACATTTTAACAGGCACTTGCGGTAATGGCTCATTTATTAATCTATCAAAATCTACTTCTTCCTCATCCAGGTAGTAAACCGACTGTCCTCCACTTGTGTTAACCTTACTAAATGATACAGCTTTATTAACTTCAGAGCCATCATAATATCCATATAAAGGTTCCACATTCAGAACACGCAGGGCCTTCGAT tpg|BK006941.2|:298267-299749 24S185= 173=7X 
 tpg|BK006934.2| 527192 + tpg|BK006934.2| 526768 - INS CCATGGACCGGTACTTTCACCTCTACGTCTACTGAGATGACTACTATCACTGGCACCAACGGTGTACCAACTGACGAAACCATCATTGTTGTCAAAACACCAACAACTGCTAGCACCATCATAACTACGACCGAACCATGGACCGGTACTTTCACATCTACATCCACAGAAATGACTACTATCACTGGCACCAACGGTGTACCAACTGACGAAACCATCATTG tpg|BK006934.2|:526308-527652 7X26=1X18=1X4=1X2=1X9=2X15=31S 220=7X 
 tpg|BK006934.2| 35864 + tpg|BK006934.2| 36227 - INS CCCCAGTGCTTCTTGACTTCATCGTATTTGTCAGCGAAGTTAGCGTCAATGGTAGAAACCAACTTAGCCAAAGCAGCTTCGTCTTCGGCTCTGACTTCAGTCAAAGCGGCAACGGCAGAGGTCTTTTGGTTAACCAAGGTACCCAATCTAGCCTTACCCTTGACAATGGCG tpg|BK006934.2|:35508-36583 62S14=16S 83S3=7X 
 tpg|BK006934.2| 210512 + tpg|BK006934.2| 210255 - INS TACTAAGAAAAGTAAAAGAAAAATATTTAAATTTAACCATTATGATTTCCACTTTGTTTTCTCTACTATATTACTTGAACAAACTCTATTTTTGGTAATGAGGGCTGGTCACAGATTACCTTTAATA tpg|BK006934.2|:209987-210780 7X5=3S 5S17=1X41=7X 
 tpg|BK006934.2| 224909 + tpg|BK006934.2| 225385 - INS ATACAAAGCACCGTCTTTGTTAATGTTAAAGATAATTTCAACACCGTTAGCGTTTTTAATTCCCAATTCCATCAACTTGGTACCCAAAGTGTATAGTTTTTCTCTGACGACTTCAGGTTCATCGTCGGACCATTCACTTTCATCGTCCTCTTCAGCATTTTCTTCTTTTGGAATTGGCTCCAAAGTCTTTTCCTCGATGTGATGGTCACCTTCGTAAACACCAATCAAGAAATCACCCTTGGCTTGTTTCAAAGTCAATTTCTTTTGTACAGGGAACGAAGTTTCAGCCAACAATACTGGGT tpg|BK006934.2|:224291-226003 7X1=1X1=1X167= 151=7X 
 tpg|BK006934.2| 439964 + tpg|BK006934.2| 440369 - INS ATCTACAACGGTATAATAAGCATAAGCATAGCCAGGGCAATTTCGTGGATGTTCGAATAGTGAAATGCAAAAGTGGCGCTGGTGGAAGTGGAGCTGTCTCCTTCTTTAGGGATGCAGGGAGGTCTATAGGTCCTCCGGATGGTGGAGATGGGGGAGCTGGTGGTAGTGTTTATATTCAAGCT tpg|BK006934.2|:439586-440747 7X142=17S 4S1=247S 
 tpg|BK006934.2| 17316 + tpg|BK006934.2| 17327 - INS AAGTAGGCAAATAGTAAGTTCAGGCAATATAGAGAAAATAATTTATTTCTACAAGTAGAGGGGCGCAGTAGAATGCATTTGTATAGCATAGCCAAGTCAACAACAATACTGCGTTTTCTAAGGCATATTTTATTGCCATTTTTGCATCTCTCTATTCATTTTACT tpg|BK006934.2|:16972-17671 7X223= 145=7X 
 tpg|BK006934.2| 466203 + tpg|BK006934.2| 465601 - INS GTTCAGAAGCACAATAATGAGTGACGCAAATGCAATTTATGACTAATTCATCACCAAAGAGAAATATGCAGCGTTAACTCTCAATCTAAGAATATGTAACAGATTTTAATCTCACGAACTAGCGACTTTAATTGTTGTACCTTATTCCTTAGTAACGTTAGTAG tpg|BK006934.2|:465259-466545 7X5=187S 82=7X 
 tpg|BK006934.2| 165418 + tpg|BK006934.2| 165831 - INS ATAGTGTGAACTATTACTATTTTCGAAATAAGCCAAATGATTGTAACCACCAATCGGAAGAATATCAACATAACCATTATGAGGCCTATCAAATGTTTCATTTGCCGGAATAAACAGAGTATTATGAGTAATCTCCCACCATCCTCCGTTAGAACTTTCGTTCCTTACCACGTTTGAAGTC tpg|BK006934.2|:165042-166207 7X48=42S 17S1=154S 
 tpg|BK006934.2| 283755 + tpg|BK006934.2| 284058 - INS GGACAGTACTGGAGTAACAGACTTTTCTCTTGAAGAAACGTCAATTTCATTTTGCAGTTTAGATGTTCGACTAGTTTTTTTCTTTTTCAAAGTGGGTGGAACGGATCCTGAGCTTGATGCAGCTCTTCTCTTTTTCACGCTACTGTTACGCACAACTGAACTTTCTCTAGAGGCTTCAGCAGCGCTATCCATGTCTCCATCTTCTTCCACGGGGGCTAGAACACCATCTTCCTCCAATAAAGCGATGTTTTTTTCCAACTTATTCAAGTGTCTAGCAATTAGAAACAAGGC tpg|BK006934.2|:283159-284654 14S267= 5S141=7X 
 tpg|BK006941.2| 906994 + tpg|BK006941.2| 907415 - INS ATATAGACAACTCCCTCCATGCAAAGAAGATTGAACAGACTGGGTATTCAAAAGACCAACCCCGATGATCTAACACCCGAAGAGATCAACAAATTCGCCAGATTGAACATTGACCCGGACACTATTACTATCAAGAGGGTGGTCGATATCAACGACAGAATGTTAAGACAAATCACCATTGGTCAAGCCCCTACCGAGAAGAACCACACAAGAGTTACTGGATTCGATATCACCGTTGCTTCTGAATTGATGGCTATTCTTGCTCTTTCAAAGGACTTGAGGGACATGAAGGAACGTATTGGAAGAGTCGTTGTTGCTGCTGACGTAAACAGGTCTCCAGTCACTGTTGAAGATGTGGGTTGTACCGGTGCCTTAACCGCTTTATTAAGAGACGCTATCAAGCCCAACTTGATGCAAACTTTAGAAGGTACTCCTGTCTTGGTCCATGCCGGCCCATTTGCCAACATCTCTATCGGTGCCTCTTCTGTTATTGCTGATCGCGTGGCTTTGAAATTGGTTGGTACCGAGCCAGAGGCAAAAACAGAAGCTGGTTATGTGGTTACTGAAGCAGGGTTCGATTTCACTATGGGTGGTGAAAGATTCTTCAACATCAAGTGCCGTTCCTCTGGATTGACAC tpg|BK006941.2|:905706-908703 7X226= 618=7X 
 tpg|BK006934.2| 522336 + tpg|BK006934.2| 523101 - INS ATGTAGCAGTGCATCGTGGGCATCTTGCGATTCCATTGGTGAGCAGCGAAGGATTTGGTGGATTACTAGCTAATAGCAATCTATTTCAAAGAATTCAAACTTGGGGGAATGCCTTGTTTACCGGAGACCAACCCTTAGTTTGAAGTGTGCGCTACCAGGGAATCTTCTTCGGTCATTATTTTCTATCTTCACGATAATCG tpg|BK006934.2|:521922-523515 7X13=280S 16S84=7X 
 tpg|BK006934.2| 161298 + tpg|BK006934.2| 161024 - INS AGTGTAATAGATTCCGCCTTATCTTGGTATTGCCCTTTGTGTAGGCTTAAGTGTCGTGGGGGCAGCATGGGGTATTTTCATTACTGGTTCATCCATGATTGGTGCCGGTGTGCGTGCTCCAAGGATTACCACCAAGAATTTAATTTCCATTATTTTCTGTGAAGTGGTTGCCATTTACGGTCTGATTATTGCCATTGTCTTTTCTTCGAAATTGACTGTGGCTACTGCTGAGAACATGTACTCGAAATCAAACCTGTACACTGGTTATTCTCTTTTCTGGGCAGGTATCACTGTCGGTGCTTCCAATTTGATTTGTGGTATCGCTGTCGGTATCACCGGTGCGACTGCTGCC tpg|BK006934.2|:160306-162016 7X8=154S 9S332=7X 
 tpg|BK006934.2| 445801 + tpg|BK006934.2| 445273 - INS GGATGAAGACGAGTATATATATGGATGTAAAATGTACTTTATGGAAGAACAAGCCACCACATGTTGAAAACTAGATAGGCAAGCAAGATTTTTCATTTGTAGAGCTCTTACGCAAGATTTTTAAACTTCCGCTTTTTTAATCCATGAGATTCCTTTGGACACCCTTTCCGGCAC tpg|BK006934.2|:444911-446163 7X194=1S 153=7X 
 tpg|BK006934.2| 121213 + tpg|BK006934.2| 121239 - INS GGTGGACGGTCCTTTCTCAAAGAATATAGTAATTGCCATACAATATTGTAAATGAAAGGAATTATTATGATCAAAGAGATTCTTTGGGCCAATGGTAAAGCCAAGAAATGACTTAAACCAATGTTTACGTATTCCAATGCCTCTCCAACGATTGACTTGGTAGCAGACATCCTTGTATTACTCGTTTGTTCTGTTTCTATTCAAGCCTGCTGCAATTG tpg|BK006934.2|:120763-121689 7X176=21S 1S1=250S 
 tpg|BK006934.2| 422305 + tpg|BK006934.2| 422780 - INS GCTGACTTGATACGCACATCGTTGACATCGCTGACTGCAATAGGAAACTGAAATAGACGGCAAACCATTAGTTCATTCGAAAGAACGTATTGTCGAGAATTATCACTCACTATATCAGAAAATTGACACACGAATTATATAAACGAAGTTATACAGAAAAAGATTAAAGAAAAGAAAAATGTCTACATCATCCGTACGTTTTGCATTTAGGCGGTTCTGGCAAAGTGAGACAGGCCCCAAGAC tpg|BK006934.2|:421805-423280 22S93= 122=7X 
 tpg|BK006934.2| 261632 + tpg|BK006934.2| 261841 - INS GAGCAGGAA tpg|BK006934.2|:261600-261873 7X3=1S 5=7X 
 tpg|BK006934.2| 57879 + tpg|BK006934.2| 57772 - INS AAGGGAATGATGCCATTGAGGCGTAAATCTATGCCCAATTCTTGGTCATCCCCTTCTTCAAAGAGTGTGAACTCTGAAAATGAAAGTGTTAATGGTGGTGATGAGAATTCCGAATTGCCTTCCGAAATTCCTGAATCATCTGGTAGATATAATGCTGCTAATTCCTTTACCACATAT tpg|BK006934.2|:57404-58247 7X54=34S 3S1=198S 
 tpg|BK006934.2| 66303 + tpg|BK006934.2| 66240 - INS TTACCTGCTGCTGTTGCTGTTGCTGTTGCTGTTGCTCCACTTTTTGTTCTTCACAGTTGGCATAATGAAACGAAGCATGATGCGGCAGTGATGTACTGTGGACGCTGTCGAACCAATTTGTGGGTAAGTTTAGAAGACTTTCCCGAACCTGAGATCTTGCGGGC tpg|BK006934.2|:65898-66645 11S74=45S 37S4=7X 
 tpg|BK006934.2| 424191 + tpg|BK006934.2| 423954 - INS CCAAAGCATATATGGTTAACAAATTATTTGGTGAAAAAACATCCTGGTTCGTTAATGAGGAAGCTTTTGGAAAAGTTCAAACGAAAACTTTTTAGAAAAGACACACATGCGAGCTTTCGAACCTCAGATGCTAATATTACGTGTTATATATACCAAACTTTATAAAATGACATAGATATTTTATGCTGTGATAGCT tpg|BK006934.2|:423548-424597 7X4=194S 184=7X 
 tpg|BK006934.2| 6650 + tpg|BK006934.2| 6464 - INS CCTTCCAAAAGACCGTTCTACCTCAAGATGTTTTCCGAAACGAATTGACCTGGTTTTGTTATGAAATTTACAAGTCTTTAGCGTTTCGCATCTGGATGCTGTTATGGCTACCACTTAGCGTCTGGTGGAAACTTTCCAGCAATTGGATTCACCCACTTATAGT tpg|BK006934.2|:6124-6990 7X5=241S 82=7X 
 tpg|BK006934.2| 80800 + tpg|BK006934.2| 81319 - INS GGATCGGCCATATCATCAAC tpg|BK006934.2|:80746-81373 7X1=1X8= 10=7X 
 tpg|BK006934.2| 515394 + tpg|BK006934.2| 515119 - INS ACAGTCTCGTCAGTATGTACCATTATCAGATTCCTCTTCAGTATGTACAGTTGTACCATTCAGTAAACTAAACGTACTGCCGATACCGCTGGCGTCTCTTAATTTAATTCTTTCCCTTTGTGAGATGCTTGCCAATTTTTGCCATTGCTCTTTGACCTCTCCTGTAGTATCCAAAAGCATGGATCCATATATA tpg|BK006934.2|:514719-515794 7X7=6S 169=7X 
 tpg|BK006934.2| 392396 + tpg|BK006934.2| 392252 - INS ATCCTATAACC tpg|BK006934.2|:392216-392432 7X3=2S 4S2=7X 
 tpg|BK006934.2| 267555 + tpg|BK006934.2| 268130 - INS CCGTCATACTCCGTGGAAATTTACTTCTAAAAGGAGAAACAGCGATCTTTGCCGCATAAAGCCAGCCACTACTGGCGTGGAAAGATTTTTAGATTAGAAGACAATACAAAGCGGCAACGTCATAACCTTGGTATTTATTGGGCAAGCATTTTCATATCAGCGTACATACACCAGCAATGGGAATGTAAAGAAGAGTCGTTA tpg|BK006934.2|:267139-268546 7X3=6S 101=7X 
 tpg|BK006934.2| 508135 + tpg|BK006934.2| 508595 - INS GAACTATAAAGC tpg|BK006934.2|:508097-508633 7X6= 2S4=7X 
 tpg|BK006934.2| 13075 + tpg|BK006934.2| 13628 - INS GTTCAATGGAAGGTGAGACAGTGATCCTTCCAAGGGACATAACCCCCAGCAAATGCGCTTATTTCTTAAAACAGAATATCGTATTCATTTCATATATTTTCATCCATATTATTATTACCATAATCTTAAACCGCCTGGCATTATCTGCACACGGTAATACTT tpg|BK006934.2|:12737-13966 7X6=14S 142=7X 
 tpg|BK006941.2| 633145 + tpg|BK006941.2| 633353 - INS GGAGTCTCCTATTATATAGACCTTCTGAGGCTATGACTATGGCTACTAATTGGGAAATAGAAAGGTAATTACTGCTCTGTAATTTTCCTATGTCAAAGCATTTGAAACTTTGGTCGGAATTGAAGGTTAACGAATCATAGCCGTGTCTACGTGTAATTTCTGTGCTGGAAGTATTGTTTTTGAGATTGGAGTCTCCTACTGTGAAATTCATGGAATAGAAGTTTTTATTGGCACTTATATTATGCTTTGTTTTCAAGTGAGATCTAAAGGTTTTTGTCAAACTTGCATCGCTTCTTGTTAGTATCTCTCCACAATGTTTACATTTAACTTTCGTTAATTTCTTTTCAATTGCTAGAAAATGGGACCAGAACTTTGCTATATTCTTCTTGAGCATTTGAACCGGAATCCATATATTTAACCCATCATTTATGATTTCGTCTTCCGGATGAATTCTACTTGATAGGATTTTATTGCCGTCTTTTTCTATAAGTTCTATATCCTCAGTATCGTCTTCTTCCTCGTCTTCCTCCTCATGACTAGTAGAG tpg|BK006941.2|:632041-634457 7X306= 5S523=7X 
 tpg|BK006941.2| 1038502 + tpg|BK006941.2| 1038581 - INS CGTTTAAGGTGTTCGCATCCATTCTTTCAGCTACTAATTTAAGAAATTGTTCTCTTCTAAGATTTGTCAATTCTACGCCCTTTGGGTCTGTAGATGGTGTATCATTCGGATATAGTGCAATATACTTTTCAGTTTTGGGAAAATTTATCACGTAACATAATTCAATTTTAGTGGCTCTCAACTTTTGTTGTAAATCTTTATCATCTGCGCCAGATTCTTTTATTTTCTTCAATAATCTGTTATATTTTCTCAATGCTTT tpg|BK006941.2|:1037970-1039113 7X3=238S 130=7X 
 tpg|BK006941.2| 294954 + tpg|BK006941.2| 294294 - INS GCAGAAGCCCTATTCCAGTCTTCGGAAAATACCTCTCGAACAATTATCTCTGGAATTTTCAGCCGTCGCCTGCGTATATAGGCCAAGGGATAATAATGGGTCTTCCAACAGTATCGTATATGCTTATCGGGTGCTTCTTAGGCTGGGGTGTGTTAGCACCATTGGCGAGATACAAAAGATGGGTACCACCAGATGCTGATGTCCACGACTGGGAGGAGGGAGTGCAAGGATGGATTCTTTGGTCGTCGCTTTCAATAATGGTTGCTGACAGTGTAGTCGCTTTTATTGTTGTGACAGTGAAGTCCATTGTGAAATTTATTCTTATAGATGACAAAGCTGCTTTACTGAACAACATAATCGATGATACATTTCAATCTATGTTACTGGAGGAGGAACGCGCCATTAATAGCAGCAGAAGAAATACATATGTTGATGGAAGGCAGGACACCGTAAGAT tpg|BK006941.2|:293368-295880 7X5=216S 442=7X 
 tpg|BK006941.2| 800613 + tpg|BK006941.2| 800544 - INS GTTTGAATTCCTAAAGATTGTAAACGCGCTTGGGAAATTTTAAATAGAATTGAAAACTTTCCCGTAAAGATAGAGCAAATAATCCCACCAAATTATAAGGACCATCTTAGAGAAACAGCAAATAAAAATTCTCAAAAGCAGGTATTACAACTTAATAGAGATTCGTACCCCTTCGAGGCGGGTTTGGAGCTACCTTTCGAAATGGTGACAGAAGTCCCCATTCCTAGGCGACCACCGCCACCACAGGCTGCAAATAACACAAACTCTGTATCAAATAACACAAACATTCAATTCCCCGACATACTAAGTAA tpg|BK006941.2|:799908-801249 7X161= 292=7X 
 tpg|BK006941.2| 877976 + tpg|BK006941.2| 877292 - INS AGGCACTGAGTACCACCGTTGGCTAAAACTGCGAAATCTTCTTGGGCTTGGTCATACCTGCCGTAAATAGAACCACCGTCAGCTTCAATAGATTCCCAAGAACCAGATTGGTCACCATATGTGTACTTTTTACCGGTAGAATAATCAGTTACAATGACCTTTTCAATGTACATAGTGAATGGAGCGTCATTGTAGTTGGTTTCACCACCAGCCCATTCAATGGTACCAGCAGCATTGTCTGGGTCACCACCGGCCCAGATACCCATCATTAGGTACATAGGAGATTGTGGGTAACCCTCACTTGATGTGTTTGATAATACTCTGACAGACTCTCCATCGAGGTACCAAGTCGTCTTGTCC tpg|BK006941.2|:876558-878710 7X6=203S 338=7X 
 tpg|BK006938.2| 461744 + tpg|BK006938.2| 461562 - INS GTCCGTACTGAAAAATAGCTGGTGGACTTCTACACAGACAAGATGAAACAATTCGGCATTAATACCTGAGAGCAGGAAGAGCAAGATAAAAGGTAGTATTTGTTGGCGATCCCCCTAGAGTCTTTTACATCTTCGGAAAACAAAAACTATTTTTTCTTTAATTTCTTTTTTTACTTTCTATTTTTAATTTATATATTTATATTAAAAAATTTAAATTATAATTATTTTTATAGCACGTGATGAAAAGGACCCTAAGAAACCATTATTATCATGACATTAACCTATAAAAATAGGCGTATCACGAGGCCCTTTCGTCTCGCGCGTTTCGGTGATGACGGTGAAAACCTCTGACACATGCAGCTCCCGGAGACGGTCACAGCTTGTCTGTAAGCGGATGCCGGGAGCAGACAAGCCCGTCAGGGCGCGTCAGCGGGTGTTGGCGGGTGTCGGGGCTGGCTTAACTATGCGGCATCAGAGCAGATTGTACTGAGAGTGCACCATAAATTCCCGTTTTAAGAGCTTGGTGAGCGCTAGGAGTCACTGCCAGGTATCGTTTGAACACGGCATTAGTCAGGGAAGTCATAACACAGTCCTTTCCCGCAATTTTCTTTTTCTATTACTCTTGGCCTCCTAACGACATTACTATATATATAATATAGGAAGCATTTAATAGACAGCATCGTAATATATGTGTACTTTGCAGTTATGACGCCAGATGGCAGTAGTGGAAGATATTCTTTATTGAAAAATAGCTTGTCACCTTACGTACAATCTTGATCCGGAGCTTTTCTTTTTTTGCCGATTAAGAATTAATTCGGTCGAAAAAAGAAAAGGAGAGGGCCAAGAGGGAGGGCATTGGTGACTATTGAGCACGTGAGTATACGTGATTAAGCACACAAAGGCAGCTTGGAGTATGTCTGTTATTAATTTCACAGGTAGTTCTGGTCCATTGGTGAAAGTTTGCGGCTTGCAGAGCACAGAGGCCGCAGAATGTGCTCTAGATTCCGATGCTGACTTGCTGGGTATTATATGTGTGCCCAATAGAAAGAGAACAATTGACCCGGTTATTGCAAGGAAAATTTCAAGTCTTGTAAAAGCATATAAAAAT tpg|BK006938.2|:459332-463974 7X7=842S 77S42=1D134=4I297=7X 
 tpg|BK006941.2| 173647 + tpg|BK006941.2| 173911 - INS CTTTTTTTTTGTAGAACGCGCTTAGAAAATGGCATAAAGAAAATGGCTATTTGACTTGATTTTGAAAGTTGTTCTCAAGACTCGAATGGTGGAAGATAACAACAGGACGTTTATTACATGGCATTGCATCAGTATTTATCAG tpg|BK006941.2|:173349-174209 7X6=65S 65S6=7X 
 tpg|BK006941.2| 580451 + tpg|BK006941.2| 580522 - INS GTACACCATGCCTCTTATAGTAACTGTATATCTTCTTAACAGAAAGAACACCGGGATCAGTTTCTGCAGTATAGTCTTTGCCTGAAAGGGCCTTGTAAAAGTCCATAATCCTTCCAACAAATGGGGAGATCAATGTGACATTTGCCTCCGCACAGGCTACTGCTTGCGTAAAGGAAAACAGTAATGTCATATTACAATGAATACCATGCTTTACTTCCAATTCTCTAGCAGCTTGGATACCCTCCCAC tpg|BK006941.2|:579941-581032 7X218= 124=7X 
 tpg|BK006941.2| 331241 + tpg|BK006941.2| 331374 - INS TTGGTCCTCAAAGATATCTTCTTGGGACATTAATATTAATGTGTTTGAAGTCATTATTCAAACCATGACCAACAAATACGCATCCGAGCTGCATTAAAAGCCAGACTTTTCGATATACAACGTTTCTTCTCACAAGCCTTTTGGTACTCTTTTCAGGGTCCAAGTCACCAGGAAGAATCCCACTATATCTTGTCAAATAGTCTTCTATGTGGTTCGTGTTTACCACATAATCATCGACAAATGGTACTCCATACAGTTCTCCTTCTTCGCCTCTAATAATGGATATTCTGGCCAAAGCAGTTCTTTTAGGTCGAATAATACTTCTGATTCCTTGATGATCGATTTCACATAGTTCACTTTGTAATGAGACAAATTCGGCATCAATGGCAACCAAGGTTCCAGATTTAGGTGCCTCATCATGTGTTAATAACTTATATTCACGTCTTGCAGTAT tpg|BK006941.2|:330321-332294 7X164= 4S435=7X 
 tpg|BK006941.2| 65511 + tpg|BK006941.2| 65701 - INS GTCTACTCTAGTGTCATGATCATGGAAGAGCTTTTGAAGCAGTGTCATGATCATCGTCATCATCATTTTCAAGTTTAATTAGTAATGCATAAAAATCTTCCATATGCATAGTGAGCTCATATAACAAATGGCCCAAATAGACTGGATCTCTTTGAGAAGGCGGATTGTCTACTATGGTGGTACTTAACAAATCTACTTCGTCATAGTCGGAATTATTCTTCCTGATCAACTCAATTATAATAGATACGGCAACTCCCATTGCATGGCCTCTTTGAAATAAGATTATATTAATAAGTTGGTCGACATATTGCGGAGAGGCAAGCTGTCTTGTCAATCGGTTAGGTCCGATCCACAAAGTATCCAGTTTAAAATTGGTGGAAATGCTGATCAGTGCTTTTAGAAGCTCTCCGCTACTGTTTTGAATACCAGGTGAGTATTTGCTATTTTCCAAGAGATTCAAACACTTAGGTATCAGA tpg|BK006941.2|:64545-66667 7X161= 7S455=7X 
 tpg|BK006941.2| 652095 + tpg|BK006941.2| 651359 - INS ATATTCAACAAGGTATGATGCGGCAGTTTCAGTTCAATTAGTCTGATCACCGAGTTTTTCTGGAACTCTGAATCAGTGGTTAAGGCATCCCACTCACCCGTAGTGGCGATCTTGTGATTTTCGTACTTTTTCGCACCAAATGCGGGCAACAGGGCGAGGTGATCCCAGGTCTGGATTTCGTTGTACTCTGCGTGAGGCCCATGAATCAGCTTTTCGATAGTGTAGCCGTCGTTGTTAAGGACAAAAAGATACGGCTTTAACCCCCATCTGA tpg|BK006941.2|:650803-652651 7X4=221S 5S250=7X 
 tpg|BK006941.2| 333593 + tpg|BK006941.2| 334348 - INS GGAATCTCATCGAAGCTAATCGCTGTAATTTCCTTATCCCTATTATCGAAGCGAAAGTATGGCTTCTTCAAATGTTCCGAAAGATCAACTGGATTGTTGAAGAAATGTTGCCAATTATTCATAATACATTCACCATTCAGAAACTCAGTATAGCAATTGTGTTCTAGGAATCTCTTAGGGTGTAATGCAGTTCAAAACAAAAAATAAGCAAATAAAAAAATTTTCAGAATGTAAAAATTCTAGTTAAAATGAACGTGTATTATATGGTAATGATGTGTCTCTTGGAGATTCTATTTCTTGTGTTCCTCTATGCCCACATAGTACGTTAT tpg|BK006941.2|:332921-335020 7X8=272S 4S161=7X 
 tpg|BK006941.2| 721023 + tpg|BK006941.2| 720785 - INS GGTCCCTCTGAGGAGAAGATGAAGGAAACGCTGCAGAATCAGAAAGTGACAACGTCGCTGCATCAAGGCAAGATTCTACGTCTAAATTGGAAGATTTCTTTTCTGAAGATGAAGAAGAAGAAGAATCTGGTTTACGCAACGGTAGGAACAATGAATATGGGCGTGATGAAGAAGACCATGAAAATAGGAACAGAACAGCTGACAAAGGTGGAATCTTGGACGAATTGGATGATTTCATTGAAGATGATGAATTTTCTGATGAGGACGACGAAACCAGACAAAGGAGGATCCAAGAAAAGAAGCTTTTAAGAGAACAATCCATCAAACAACCTACACAGATTACTGGTCTATCGTCGGATAAGATTGACGAGATGTATGACATTTTTGGTGATGGTCATGAC tpg|BK006941.2|:719969-721839 7X170= 4S385=7X 
 tpg|BK006941.2| 792113 + tpg|BK006941.2| 792764 - INS GCCCAATTACATCTGCCCATGTACATGTTTATATTTATCTATCTGTTAGGACTTGTGAAACAATGCTATTTTCCTGTGCACTATGGACTATGGCTTTGCGTTTACATTTTATGCCTCCAATTTTTCACAATCCTGTCCGACGCTCAGATATTGGTGTGGAAGTAGAGCTAACTCTCTATCTCAGAAAAAAGGTTAGAGCAAGGCAGATCTTTTGCAATAAGAATCAGTTACCATCGATCGATTTGAATTCATATTACTAGTACTTTGCAATACACTGTGTAAGAAGATGTCATAAAGATTGAGAAACGGTCATCAAACTTAATGTAAGCAGAGACACGAGGATTGATGAGGAAGTAAGATAATGTGCGACAAGGAAGAAAAAATAATAGCATTATGT tpg|BK006941.2|:791305-793572 7X86=1X393=2S 75=1X249=1X47=7X 
 tpg|BK006941.2| 1072023 + tpg|BK006941.2| 1072532 - INS AGTATTTTACAGAGAAGATAGATAAATGCCAGTTAATTTTAGGAGGCAAGATATTATTGTCATTTATGTTTGCCATTTAAAGCAACATTTTTATGGCAGAACATAACATTAAAAGAATCCGATCTAAATTTAACTATAATAGTTACTAGATACGGACATATCTCTAGGAACTATGAAGGCTGAAATGTCTAGAACTTTGGAAAAGAGATGTCCTTTCTGCGTAGCTTAATTCATTTCCTTCCTAAAAAGTCCGTAGAAAGAACACTGCACCTCGC tpg|BK006941.2|:1071459-1073096 7X189= 138=7X 
 tpg|BK006938.2| 28766 + tpg|BK006938.2| 29033 - INS TCAGAGAGGAGTTGGAAATGGGACAATGAGATATACCACAGCGACGCTGTTTAATCACACGCGCTTCGGCATCTGTTAGATGAATACAATGTGCCAATACTGTTTTTTCTGTGAGCAGCCCATATTTGTCGTATACATCAGTATAGCTCTCACATTCGGGAAATAAATCTTGAACCC tpg|BK006938.2|:28398-29401 7X6=82S 85S4=7X 
 tpg|BK006941.2| 531407 + tpg|BK006941.2| 531115 - INS CCAAGTGCATATACATATATACTTAATATTATAAACGCATATACTTTTATAAACTTGGAATAAGTATTATATATTTATTTTGACCATCCGGAAATGCTTTATTTTACACTTGGAAAGAAAAGTGCATTTGGAAAACTTTTACATGTCACCCAAGTGCATACTGCTGACGATACAGGTTTAGAGACTAAAGAGAGCGCATGGAAGAAAACTTCAAAGGAAGAGAAGAAGGATCGCAGAGTTCAAAGGAACTCTTAATTTGGGCC tpg|BK006941.2|:530575-531947 7X5=179S 247=7X 
 tpg|BK006938.2| 1476445 + tpg|BK006938.2| 1476699 - INS GATCTCAACCAACCACACACACAAACACTAATTCACTCTCACTCTCTCACTTTCCCTTTCGACGACACACACAAAAAGACTTTCTGGATGCCCCGCGTTTTTTGTCACTTGATTCTTCGAACAAAGACGCAGGCAACTACCCCTGAAGGGCCCACCCGAAAGTAGTTGCTACTGCTCGTTGCGGTGGCTGCCAGAGTGGCGACGTAGCGTTGCGTTGTGGCTAACATTGGTGAGACAACCCGATTAAATTACTTAATGGGCTCTCCCACCGCCTTTGCACCCAGTGACAGCCATTTTGAAGATAGCATCGGGC tpg|BK006938.2|:1475805-1477339 7X5=223S 294=7X 
 tpg|BK006941.2| 599383 + tpg|BK006941.2| 599540 - INS GATTGCCACCAGCCGCATCTTACAATGTATGCCACGATACCGCCAGGCAATAAATGAATATGGAGTGTCACTTCGGCTCCGTAAGCCGGCGCTGCATCCGCCACCACAGTTTTTTTTAGCGTCGCTGTCGCCGCTTTGCCACAGAAAAAGAAAAA tpg|BK006941.2|:599059-599864 7X4=73S 72S6=7X 
 tpg|BK006941.2| 579891 + tpg|BK006941.2| 579667 - INS GGACAATGCCACCAGAAGGTTTTGATATTGAAGAACATAGGATTTTTAGTCAGTTTTTGGTGATTATTTCAAATATTATTGAGGAGTACGATAGAGATATTCAAGTGGCAGCAACGCATGTTAGGGCATATCCTTCAAATTTGTCGGTGCAAAAACAACGCCCTCTTATCTCAGACAATGCACCAAGTTTGAATCATATCTCAACTGCGAGAGAAGTTCATTCGAACATAAAAGTCACAACTCCCAATCGCAAGCAGACAGAGGACAATGCCACCAAGGGAGGATTCAACATCAGCAAACTTACTCTGAAGGTCAATAAGCCTTTCAAGAAGCCCAAGAGGATATTAAGTACTAATGTGGTAAATGAATCAAATAGACCGAGCATAAGG tpg|BK006941.2|:578875-580683 7X192= 365=7X 
 tpg|BK006941.2| 277755 + tpg|BK006941.2| 278382 - INS TTTTTTTTTTTTTTTTTTTTTTTTAAAATCTAAATATGTTGCTTGAATTATAAATACAATAACGGGAAAACATATGATGTGTCATGTTCAAAAAGCTTTGAATAGGTGTCTTCCATCAAAAGGGTCACAGGAACATGAATTTCGTTCCGTGATTTTAATAGTAATCAGTTCATTTCCGTATCTTGTTCTTGGTGCGTAAAACTGGTTTGCGGAGGAGCATTTTCAATTATTGCGTTTTCTGGCAATGCAAATGGCCTTTCATTGGTAGGAACGTTTGAATTGGGTGCAGCGC tpg|BK006941.2|:277157-278980 7X199=20S 1S1=189S 
 tpg|BK006941.2| 684418 + tpg|BK006941.2| 684252 - INS AAATGCCTTATTGGCTTTTCCCAAAGTTATATTTTGAAGACAGGTTTGCTCTGTAATCATATAGTATCTGTGAAGAAAATGCAGACATCTGTAGACGATAATAGGTTCCTCTAAGTCAGAAATAATTCTAGACAGTTCTTTACTGTAGAACTCACAGTCTCTGGCAGAACCAATGCGTATATGTATTTTAATGAGTTGGAAAAAACTAAACGATAGACTTTTTAGTAATGCTAGCCTGGAT tpg|BK006941.2|:683756-684914 7X147=33S 4S1=216S 
 tpg|BK006941.2| 773350 + tpg|BK006941.2| 774007 - INS CCCTTAGCATGGGAGGTATACTGGAATATTACGGCTCTTTTTTTTTAGAAACATATTCCTCAAATGGGTAAACGGACCCTGGTGCAAGGTGTGGGTGCTGAGACAAATACGATCTGAGTTGTTTTAAAAAGGAAAACAAATGAATGCGTGCCCAAAGCGGAAAATTGGTCAACATCGATGCGTAATTAGTAGGCCCAGGTGAGCCTGTGCCGAACATGTATCTCTGCGCAGATTACTATATATTCCCGAGCATAACAGCATATAGTTTTCTGTCACATAGGCCTTCCTCCAACTGCCATCACTGTACATAGA tpg|BK006941.2|:772712-774645 19S144= 62=101S 
 tpg|BK006941.2| 393857 + tpg|BK006941.2| 394022 - INS GTTGATGACATCCTAGCATCCATATTGACATCCATTCAAAGTTTATTCAACGATCCAAATCCAGCTTCGCCAGCAAACGTTGAAGCTGCAACATTATTCAAAGATCATAAATCACAGTACGTCAAAAGAGTTAAGGAGACGGTAGAGAAATCTTGGGAGGATGATATGGACGATATGGACGATGATGATGATGATGATGACGACGACGACGACGACGAAGCAGACTGAGAA tpg|BK006941.2|:393381-394498 22S100= 107=16S 
 tpg|BK006941.2| 751477 + tpg|BK006941.2| 751081 - INS GTTTTACTTCCTCAGTATGATATTCATACAAGGAATCGTCCTTTGGAAGGACGCTCGTATTCTTTTGTGAACGGTCATTTGGTATTTTGTGGTTTTCAGCCGCGTGTATACCTTCAGCTTGTTTGTGCTGCCTACTCAATATTTCTTGCTTCAAGGCCTCATCAGCGTTTTTCTGGCGAGTTTGTTCCTCGATAGCCTTTTCAGCTTGTAATCGCGTTCTTTCCCTCTTGACTGCCTCCAGTTCTTTCTCTTCGGTTGCCAGCTTATCCTGTAGTTCAGTCAATTGGTCATTATAGGTTTGCTTGACT tpg|BK006941.2|:750451-752107 7X316= 154=7X 
 tpg|BK006941.2| 90041 + tpg|BK006941.2| 90746 - INS GTACTCCATATGGACCTCTTAGGTGAGTGATCTTATTAAAAAAAATAAAAAAAATAAAAAAATATGAAAAAAAAAGAAAATTAAAAACTAAACAAATTTTATGACAGGAATAAAAACTATAAAAAATGAAAACCAAAAAAAAAAA tpg|BK006941.2|:89737-91050 7X5=67S 66S7=7X 
 tpg|BK006941.2| 612198 + tpg|BK006941.2| 612318 - INS GACCGTATCCATCACCATAAGAGAAACCACCACATGCGGCAAGACCGATGAAGTCATCCAAATGGAACCTACCTTCTAGCAAATCTGTCATAGTGACATCCACTGAGTTGAATCCAGCTTGTTGGAAGCACCATGCCATTTCCATTTGACCGTTCACACCTTGCTCTCTTAAGATAGCAACCTTTGGCCTTTGACTGGATAATTCTAATC tpg|BK006941.2|:611764-612752 7X188= 197=7X 
 tpg|BK006941.2| 428800 + tpg|BK006941.2| 429353 - INS GGGTAGATATAGCGGGGACTCAAAGTTTAGCATCCACTTTAAATATCATTCAGTTCCTTCTATCGAAATTCTTAATCAACATGGGCAGTATTTCGCAATTAATTAATCAATACAACAGGAAATGCATCACTACTAATAACATCAATAATAACAACATTAACAACAATGGCGTTATTAATGGTAGTACTAACACCACTAGTACTACTACTACTACC tpg|BK006941.2|:428356-429797 24S90= 96=19S 
 tpg|BK006941.2| 390882 + tpg|BK006941.2| 391383 - INS GGCTATGTTTTTCTGCCGCCAAGCAAAAGAAAAGAACGCAAGGTGATTTACTCTTGGTACTAACATATATGAAATTTTTTGTTAGTTTAAGGAACAAATGGGATTTGGGTCTGTTAACACTCATCAATAAAGAAATCTCCGAATCATTTCAAGGAGAAGGTGAGCCTGAATTAGCATTCATCAACATTTCCAATAATACTC tpg|BK006941.2|:390466-391799 10S45=52S 96S5=7X 
 tpg|BK006941.2| 871866 + tpg|BK006941.2| 871919 - INS GCTCTACCTGAAGCTTGATTGGAAGCTTGACCGCTATTTAACAGTAAATCAAATATAACGCCCCATATTTCTTTTTTCCAATACCTTTTGAATGGGTTCTTCAATTTGCATCGTCCATTCTGCAGCTGGATTGTTTCTATGAATTTTCCAAAAAGCATCGAATGTATGACGCCTGCTAATCCATAATAATCCGCTTCATAACTCCATGGCTTGCCCGCACGCATTTCCCAGCAATCTTGCTGATCAGCCTTCCAATTTGATTTGAATTTCGTTCCAGGTGGTAACAG tpg|BK006941.2|:871278-872507 7X199= 270=7X 
 tpg|BK006941.2| 247113 + tpg|BK006941.2| 247291 - INS ATTATCTACTGTTACTGTTCAATGTTCAATGCCCTATCTGGACACTATGAAACCAGAAGGTACTGTTAATAGATCAGTAGCGAACGAGTTGCTTGCGTTGGGCAATGTGGCAAAAGACCATGACGACAATTCAGATTACGAATCAAATGATACTGGTGTGAATGATGAGCTAAAGCAAGCACAGGATGAAACCACTCCCACAACCGTAACATCAAGTGATGATAACAAGCCTACGTTTTCAGAGAAAATATTAAGTAAATTCTCTAGGCC tpg|BK006941.2|:246559-247845 7X233= 15S229=7X 
 tpg|BK006938.2| 837069 + tpg|BK006938.2| 837145 - INS GGTGGTAGGCATGGTTGAGATCATCGAGAAGACTGAAGTTAACTCTGGGTTCTTTTACAGTTCTGCGGACCAAAGGGACAAGTTGGCCGCTAGTGAGAGGAAGTTTGTGGATGCCAAGTTGAAGAAGATCATCGACTTGAAAAACGAAGTTTGTGGCATGGATCCAGACAAGGGTTTTGTTATCATTAACCAAAAAGGCATTGACCCCATGTCTTTAGACGTGTTTGCCAAACACAACATCTTGGCTTTGAGAAGGGCCAAGAGACGTAACATGGAAAGATTGCAATTGGTCACTGGCGGTGAAGCTCAGAACTCTGTGGAAGACTTGTCGCCTCAGATTCTTGGGTTTTCTGGCTTGGTCTACCAAGAAACCATAGGCGAGGAAAAATTCACATACGTTACAGAGAACACTGACCCCAAGTCTTGCACCATCTTAATCAAGGGCTCCACTCATTATGCCCTCGCTCAAACAAAGGATGCGGTGAGAGATGGTCTCAGAGC tpg|BK006938.2|:836053-838161 7X375= 9S477=7X 
 tpg|BK006940.2| 148628 + tpg|BK006940.2| 148503 - INS AAAGAATATCTTCCACTACTGCCATCTGGCGTCATAACTGCAAAGTACACATATATTACGATGCTGTCTATTAAATGCTTCCTATATTATATATATAGTAATGTCGTTAGGAGGCCAAGAGTAATAGAAAAAGAAAATTGCGGGAAAGGACTGTGTTATGACTTCCCTGACTAATGCCGTGTTCAAACGATACCTGGCAGTGACTCCTAGCGCTCACCAAGCTCTTAAAACGGGAATTTATGGTGCACTCTCAGTACAATCTGCTCTGATGCCGCATAGTTAAGCCAGCCCCGACACCCGCCAACACCCGCTGACGCGCCCTGACGGGCTTGTCTGCTCCCGGCATCCGCTTACAGACAAGCTGTGACCGTCTCCGGGAGCTGCATGTGTCAGAGGTTTTCACCGTCATCACCGAAACGCGCGAGACGAAAGGGCCTCGTGATACGCCTATTTTTATAGGTTAATGTCATGATAATAATGGTTTCTTAGGGTCCTTTTCATCACGTGCTATAAAAATAATTATAATTTAAATTTTTTAATATAAATATATAAATTAAAAATAGAAAGTAAAAAAAGAAATTAAAGAAAAAATAGTTTTTGTTTTCCGAAGATGTAAAAGACTCTAGGGGGATCGCCAACAAATACTACCTTTTATCTTGCTCTTCCTGCTCTCAGGTATTAATGCCGAATTGTTTCATCTTGTCTGTGTAGAAGACCACACACGAAAATCCTGTGATTTTACATTTTACTTATCGTTAATCGAATGTATATCTATTTAATCTGCTTTTCTTGTCTAATAAATATATATGTAAAGTACGCTTTTTGTTGAAATTTTTTAAACCTTTGTTTATTTTTTTTTCTTCATTCCGTAACTCTTCTACCTTCTTTATTTACTTTCTAAAATCCAAATACAAAACATAAAAATAAATAAACACAGAGTAAATTCCCAAATTATTCCATCATTAAAAGATACGAGGCGCGTGTAAGT tpg|BK006940.2|:146513-150618 7X8=486S 124=377S 
 tpg|BK006941.2| 606788 + tpg|BK006941.2| 607463 - INS GATATCAAAAACTTACCACGTCAACGTGAGTTGTTGAATGCCAAAAATGGAATTGATTTTACGCTGATGGTGGCGGGTCAAAGTGGATTGGGTAAAACCACGTTTATCAATTCCTTATTTTCTACTTCTTTAATTGATGATGACATCAAAGAAAACAAACCTATTATTCGTTATAAAAGCATTGTAGAAGGAGATGGAACACACCTTAATTTCAACGTCATCGATACACCTGGTTTTGGTAACAATATGGATAATGCATTTACGTGGAGGACAATGGTTAACTATATTGATGAAGAAATAAGAT tpg|BK006941.2|:606166-608085 7X1=1X251=22S 14S1=259S 
 tpg|BK006941.2| 556016 + tpg|BK006941.2| 556210 - INS TTTGCAACATAGATTTAAGTGTGGATGAAAATTATGTGCTCATTGTGAAAAAAAAGTTTTGCTTTTACTAACAAATTTTTTTATTATTTGTTTTCAATAGACGTTTCCTCTGACAGAAGAAAGGCCAGAAAGGCTTATTTCACTGCTCCATCCTCTGAACGTCGTGTTTTGTTATCTGCTCCATTATCCAAGGAATTGAGAGCTCAATATGGTATCAAGGCTTTGCCAATCAGAAGAGACGATGAAGTCTTGGTTGTTCGTGGTTCCAAGAAGGGTCAAGAAGGTAAGATTTCATCTGTTTACAGATTGAAGTTTGCTGTTCAAGTTGACAAGGTCACCAAGGAAAAGGTCAACGGTGCTTCCGTTCCAATTAACT tpg|BK006941.2|:555250-556976 7X3=1I118= 188=7X 
 tpg|BK006938.2| 835278 + tpg|BK006938.2| 836033 - INS CTTTCTGGAAAGCGAGGGAGAGTGAGAGGTGTGGGTTCTGCGGCAGAATGGATACGGGCCGTGGATCACTGTTTACGGGAGTTTTGCTTTGGTGGCAAAATTTTCGCTCGGTGATGTGTTAGTAGTTGTTATTCTGGTAAGAAACGAACGAAAGACGGAAAGGATTATGTATAACAGTGTATGTGTGCAGTGTGTGGAAAAGGTAAAGGTTAAGGGTGTGGAAGCAGTGAGAAGCAGAAGATTATAATATAAGTAGAGTAGAAGCATGTCATTGCAATTGTTGAATCCGAAGGCTGAATCGTTGAGAAGGGATGCGGCTTTGAAGGTTAACGTCACATCTGCTGAGGGCTTACAATCCGTCCTAGAGACCAACTTGGGCCCTAAGGG tpg|BK006938.2|:834490-836821 7X483=1X184= 6S369=7X 
 tpg|BK006941.2| 22892 + tpg|BK006941.2| 23319 - INS CCCCAGAGTACAGCTTGAAAAAAAGTGCGGGGCTCCAGAGCTCCACATTGGTGACCCCAGAGTATACTGCTCTTTCTAATGCCTTTTCCATCATGTTACTACGAGTTTTCTGAACCTCCTCGCACATTGGTACCTAGAAATGGCTATCATGCCGGACGGCACCGGGCAATAAACCGGACGGCACAAAAAAATCGAAGAAAAGAGATTTCTTTTTCTCGCGGGCAGTTTTTCCGGTCGATCGACATTCGTACGGTACTTTCTCTGTTTCAGGGACATCATGTTGTAAAAGAAAAAGACAGTTTAGGTAATCGTTCTTTTCTTTCTGAAAAATTTTCCACGACGACGACGACGACCACGAAACACCTTTGATTGCGAGATCCACGAAATTACCTCCTGCTGAGGCGAGCTTGCAAATATCGTGTCCAATTCCGTGATGTCTCTTTGTTGCACCTTCGCCACTGTCTTATCT tpg|BK006941.2|:21940-24271 7X432= 455=7X 
 tpg|BK006941.2| 415664 + tpg|BK006941.2| 416116 - INS AATATACGTTTTTTTTTGTATTTTTGCCTCCCTAGTTTCAAAATGCACCAAATTCTCCCCTTAATGCTTTTTGTTTTAAGTCCCAAATAGCCATCCTTTCATCATCGGGCAAGATAGAAATTTGACTGTCATTCAGTTGTAACACCTGTTTCAGTAGTTCTTTCTGTTTGTTAAGCACAGCTGGATCCACCACCTCGTTCACGCTATTGTTATTCGTAGCCGATGCCTCTTCTTGCGGCCTGGAAGCTAACGGGATCAAATCATCCACTTTACATATCCCATTCG tpg|BK006941.2|:415080-416700 7X162=1X64= 268=7X 
 tpg|BK006938.2| 600544 + tpg|BK006938.2| 599779 - INS GGTCAAAGAAAAGTTAAATTTTACCTATTTAGGATTTTAATCTGTTGGAGTTAAGGTGAATACGTTTTTCCATATTGGGGTATGCAGCTCGAACCTAAAGTGGTATGTACACATCCCCTCAAGCACACCCATTACCCTTATAGGATTAATGTAAGCAACAGCTTACACGGAATTGGAAATACTATTCAACGATCCATGCATCTGCCAGATTCGGACAGGCATATTCCCCAATTGGATATAGAAAATTAACGTAAGGCAGTATCTTTTCACAATGTACTTGCAACGCGGCGACTTAAAGTTGAAGTACAACCTGCAGCAGCGGCTTTTTGTACGGTACGCCAAACTGTCAATGGATAATATTGCGTAGACCGAAAAAGGTAATCCTCAACACTACCCGTG tpg|BK006938.2|:598967-601356 7X5=378S 18=1X181=7X 
 tpg|BK006941.2| 383405 + tpg|BK006941.2| 383221 - INS ATCTTGAGACATCTTTAATCTGATCTGAAGAAGTATTTCTACTCATCACTAATATCTATTCCGCTATTATTATAGTTGTAATTTATGATTCCGTGGTAAGTGATTTGAACTTTTGCTTCCTTTCGAAAATTTCAAGAATATGGTTTGGTTGTGCTGTGCAAGAGCGGTTGTATTGCGAAATAGAACCCATCGAGAAAAGAAAATGAAAAAGACGGCATTAAAGACTAGCTCTGTTTTAAGACAAATATTTACAGGCCAGAGAATAAAGAGATACTCGTATGTATGAATTGTAGCCCCTTACACACATATGTATATATATCGATGTGAACATAGCATTTATTAACAGTTCTGCTCAGTACAAATGGTAGTAGTACTAGTGATGAGGTTACTCCGACACCGTTAACAGCGGTAGTAAAGAGAAGGCCGAGTAAACAT tpg|BK006941.2|:382337-384289 7X5=207S 422=7X 
 tpg|BK006941.2| 109266 + tpg|BK006941.2| 109940 - INS CACTGAAAACCTATTACGACAAGTTAAACTCTCGTGATTCACATATTTCCGATGAAATTACAAAGGAATCTATGTGGAATGTTTATAAGTTATTTTCCTTGTATTTTATTGACAAGCATTCCGGAGAATTCCAACAATTCAAGATCTTCACTCCTGATCAGATCTCTAAAGTTGTGCAGCCACAACTATTGGCTCTTTTGCCAATTGTGAGGAAAGACTGTATAGGTCTGACAGACTCCTTTGAATTACCTGACGCGATGTTAAATTCTCCTATAGGTTACTTTGATGGCGATATC tpg|BK006941.2|:108660-110546 69S131= 148=7X 
 tpg|BK006938.2| 61783 + tpg|BK006938.2| 62516 - INS CCAGCACCTTCATCGAACCTCAGTTTCGCGAGATGAGAACCGTTTCTATGTATGGGGAAAAACCTCCGGTACTCTTCGAAATAGCGTGAAATTGCGGATTCGCCAATTCTCTTGAACGCTCGTTGGTAGAACAATCTTAAATGTTCGCACTGTGAAGGCGAGGCGATGCTGCTTATTTGGGAATGCGGGACCGGCTCACATTCGCGCACAATGGCATTCAATTTGCCGTTGTACATTTTCACTTTTATATTCATCTTACAAACTATGCCGTATTGCGAAAGGTTTTCATCGCGGCCGTTCTGTAGATCTCTTAGCC tpg|BK006938.2|:61137-63162 14S245=24S 35S5=7X 
 tpg|BK006938.2| 543967 + tpg|BK006938.2| 543929 - INS CAAACACCCTGACCGCTTATTTTCCGCGAAGTTCGTATATTTTAGTTTTCTTTTACTCCAAGGGTTCGTGACGTCGAATTCCTATCAGCTTTTTTTTGCGCTTGGCGTTCTAGGTCCCTGTGCCCGTCTGAAACTATTCGTACATAGCATTACTAGAGTACATAATATCGTCTACCATACATACGACGGGTAGCCAGATTTTGTGCCGGATTGTCGGGGAAAAGACGGCAAATGAGCTCATACGTAA tpg|BK006938.2|:543421-544475 23S107= 113=18S 
 tpg|BK006941.2| 925939 + tpg|BK006941.2| 926039 - INS GGACCGACCATTTAGGATCATATCGCCGGGAGAAGAGACAAAATATCAACGAAGTTCGTTGAGTACTTCCCTGACGAAACCTTATGGGGCAAAGGAAAATCAGAGGCCTTTTGGCACCCCAAGAGCCTTTGCGAGATCATCGTGGAATAGAATAGATCTGGTATCTTCTGTCAGTTTTTGGCTAGGTATGTTTTTATCCATAAAAAGTTATGATACAAAAACAGGCATAAGAATATTCAAGCCCCTTGCTATATTAAGGATTCTTCGACTTGTAAACGTGGATACTGGTATGCCCTCAATTCTAAGG tpg|BK006941.2|:925311-926667 7X7=183S 154=7X 
 tpg|BK006938.2| 953348 + tpg|BK006938.2| 953556 - INS TGGTGGTGTATTGGGACCCCGTTCTGTATGAACAAAAACATATGGTTTGGGAACATAGAGAACAAGATGCGTTAGAGGCATTATATGAAAACGAACCGTGGATTCGTTCGAGAATAGGATTTTTGCCCTTAAGAACGATCAATGCATTCCCACCGGGAGCATGCTCTGAATACAGTGGTGACTCAAGATACTTTTACAGTGAGAAAGACCATGATCTTGTTGTGAATATGGCCGGATGCAATTTTGGCAGAGATTGCTGGGGCGAGATGCAGTACTACACCACTTTAATGG tpg|BK006938.2|:952752-954152 41S169= 197=1X75=7X 
 tpg|BK006938.2| 1410183 + tpg|BK006938.2| 1410358 - INS CGAATAGTATCTTCGAGGGCGTGAGTCAGGAACTCGGCAACAATGATGAGTCGCAGCACAAGATCACTATCCAGCCACGCCTCTAAGGTGGAGCCCACAGGATTAGGGACCAGGAAAAAGATAGCGTGCAGTGCAGGACGATAGAGGTAGCACAATGGCGGTAGCGCCACGCCTACCAGGATCAACAAGTCTACTAGAGTGCAGGGGTACTCAACAGTGTCGATCTGGATGAGCGACAGCTTCCTCTTCTCCGCAGCGATGCGGAACATCTTGTTGAAGATTTGCTTGATTCCGGTAGC tpg|BK006938.2|:1409571-1410970 12S167= 281=7X 
 tpg|BK006941.2| 508782 + tpg|BK006941.2| 509556 - INS ATATTACATAGCATTAAATCTAAGTTTCCTTCTACGTTATTCAATTGTTCACTTTGATGACCCAGCATACCCAATGTGTTCATACCTGCTCTTTCGGCGTCTTGAGCCATTTTTAGTGTATTTCTAGTAGAGGCTACGGAACTCTGTTTCGTAAATTTGATCTCCTGCTTGATTTCATCTACTGCTTCATCTTCTTCCTGCTGCTGGCGAGCCTCCTCTTCTTTTTGTATTTCTTCAAATGTTTTGTAACCCCTTTGATCTCCATATTGGTTATTTGTTGCGTTAAAGTGTTGCTGTTGCTGTTGCTGCTCATCCATGAACCACTGTTGCTGCTGCTGCTGTCTTGAACTATGATCAACTTCGGACGCATTTAAATCTATTGAATCTTCATTCGTCATTACTG tpg|BK006941.2|:507962-510376 7X215= 378=7X 
 tpg|BK006941.2| 779040 + tpg|BK006941.2| 779504 - INS TTCCTATACCTATTATTCTATCAGGGAAATGCATCAGATAATGGATAAAATGGAAAGAATGGAAAGGAATTGTAACATGCCTATATATGGAAAACGAGCTTTTAGAGCTTTCAAGTTAACCCCGGGCGGTTAGTGTAGTGGTTATCATCCCACCCTTCCAAGGTGGGGACACGGGTTCGATTCTCGTACCGCTCAAGATTACTTTTTTAATTTTCATACTTTTTCTCCTAATATCTTGCAAATCATGACTGAATTGACATTAACTGATGCAAATGGGTGGGAAAAATGCTTATCAACCCCCTAAAAAGTCAACTTCTTCGTTAGTGATTGCTATATGTGGCGTCAAGAATTACAAGAAGCTGGCGAGCTTTCCAAGCCCCTTCAGGATTAACCGTTTTTTACCCTTTTTTTACAAATTTACGGCGGGGAATAATTCTGATACTTTCTCTTTATGAGCATTCCTCAAC tpg|BK006941.2|:778092-780452 7X141= 453=7X 
 tpg|BK006938.2| 391115 + tpg|BK006938.2| 391203 - INS TTGAGTGTGATGTTTAGTATTTCCTCTCCAATTTGCGCTTTAATTCTTTTACTTTCACTGGTAATGAAAATATAAATACTGAGGTAGACTGCAAATATGAAAATAATAATGAAATATCTGGGACCCCAGCTTAAAACAATTTTATACCAGTACGGCTTGGGTGGTAAATAGCACCATGCACTCCAAGGTTTGTAGCCACCTTGCCTGGGAGAATCGGGAAAGTTGTAGTTATTATTATCCAGTATAATAGTGGTGTCAGAATCGTCATTGAGTTTATTATAATTAATGAAGGCTAAGCTTGCTAAAATGGCAGGTACTAATGCAGTAATTGGCCAGATATATGACCTTTTTTTGTACAAGCCACCCTCCATATT tpg|BK006938.2|:390353-391965 7X268= 1S350=7X 
 tpg|BK006941.2| 946251 + tpg|BK006941.2| 946345 - INS GGAATTCCATGCTTTCACATACCCTTTTCTGGAATAGCGCTTATTTTTTCATTATGAAAAATACTAACAAATATTTTCTACAGGTATTTCTCTGAATGAACATGCAAACCTGCTTGCAGTCGGCGGCAATGATAATTCTTGTAGCTTATGGGATATTTCCGACTTGGATAAACCTATTAAAAAGTTTGTTCTTCCACATAAAGCGGCTGTGAAGGCCATTGCCTTTTGTCCTTGGTCGAAGTCTTTGTTGGCTACGGGTGGTGGAAGCAAAGACAGATGTATTAAGTTTTGGCATACATCGACAGGCACATTGTTGGATGAGATTTGCACCTCGGGACAGGTGACGTCTTTGATATGGTCGTTGAGACATAAACAGATTGTTGCTACTTTTGGATTCGGTGATACCAAGAATCCTGTATTAATAACACTATACTCATATCCAAAATTATCAAAACTACTCGAAGTTAGGTCGCCCAACCCTTTGCGTGTACTGAGCGCAGTAATCTCTCCAAGTTCCATGGCAATTTGCGTTGCCACTAAC tpg|BK006941.2|:945155-947441 7X254= 16=1X508=7X 
 tpg|BK006938.2| 575006 + tpg|BK006938.2| 575613 - INS GTATATAATAGTGAAAGTTCAGCCGCATATCTAAACCTCGATAATTTGACATACGTATATAATAGTACATGTACATAAAAAGCTACGCAAATATCGTATATCTGTTATACTACAAAACAATTACTTCTATATCATAGCCAGTTAGCGGGAACGACTTCAGCTAAATGGACTATCCATGCTTTAGGCAGAGGCGAAGCGCGGTGATTGGGTGTAACATCATCTCCTTTTCTCTACGACAAATTCCCAAAAAAAAAATTTATGCTATGTTAATACCTGCACAATTCAACCGTGCTGAAACGTAAAATTAAGGTGATTATACGGATAGTATACGATATTATCAATCTCATAAGAAAAATCTCTTTTGAATTTAACGGAGGGATTATTCATTAGAAAGCGTTCTTACCATTCACTAGGAGCGAATCCGTGGAAGGTGTTTTAACGTTGCCACGAAAAACAGCTCTACATCGAAATAAAAGACAACAATCAGTGCCCGTAAGTTTCATTACTAT tpg|BK006938.2|:573974-576645 7X206= 10S476=7X 
 tpg|BK006941.2| 154007 + tpg|BK006941.2| 154639 - INS GATACTTTCGATACCGCAGCAAAGACGAACCAAATCTTCAGGAAAATCTCTCTCTTTCCTTAATTCGGGATCAATGGAAGCATGGGACATTTTGCAAGGCATAGATAGAAGCGAATTTACACACCCGAAAGATACCGTCACAGCCCATATACTC tpg|BK006941.2|:153685-154961 8X3=1X123=11S 5S1=374S 
 tpg|BK006941.2| 151306 + tpg|BK006941.2| 151732 - INS CAATTGGGCATATATATGCATTGACGAAGCTGTATTTATCACTTGATGAAATGTACAGTAGTAAAAATGCTGTCAGGACGGGTACGGATAAGTAAGTTTCCACTTTAATGACTTGTTTGATACCGAAAATGGCAACTAAAAAGGAGCATACGGTCACTATGACAATCCCTACCCATAGGGGTACTTTATCA tpg|BK006941.2|:150910-152128 21S81= 32=71S 
 tpg|BK006938.2| 695447 + tpg|BK006938.2| 695743 - INS GATGATTATCACGTAAATACTGCCTTCTCAATGGGCAGAGGTAACCAGCAGGATGATGGCAATAGTGAAAGCAACAGCATGCATACACAACCAAGCACTATGGCGCCCGCTACGCTGAGAATGATGGGAAAAAGTCCACAGCAGCAGCAGCAGCAGAACACACCGCTAATGCCCCCGGCGGATATCAAATACGCCAATAATGGTAACTCACATCAAG tpg|BK006938.2|:694999-696191 7X4=104S 103S6=7X 
 tpg|BK006941.2| 488428 + tpg|BK006941.2| 488681 - INS TATTGCCAGACAAACCAAATCAATGTGGATAACCGCGGTACTGTGTGGTATGTTGTCTCTAATCATGGGGGTGCTAGTGAGAATCTGCCCCGATGAAGTAGCAGTGAAGGTATTTCCGGCTGCTTTCGTTCAAAGATTCAAGTACGTATTTGGACTCGAGTTCCTCAGAAAAAACCATACTGGAAAACACGACGATGAAGAAGCGCTGTTGGAGGAATCTGATAGTCCAGAGT tpg|BK006941.2|:487948-489161 7X5=111S 110S7=7X 
 tpg|BK006940.2| 270158 + tpg|BK006940.2| 269893 - INS ATCTAACAATATTCGTGAAGGATATGTCAAAATTGGATACGCTTATGTTTATGATATATCATTTATATTAATATATAGTATGCTCACATTTTCTTATTGCTGAATAGTTCTTTTTTACGTTTAGCTGAGTTTAACGGTGATTATTAGGTGGATTTTATATTAGTCTACATAAAAATAAGTGGTGGATATCTACATAAAATTGTCATAACGCGTAAACTAAAAATTATTTTTATGATCATTGAGGATCTATAATCAACTATAGACATTAATGTATGGATAATCATGAGGATTATAGGTAAATGGCAAGGGTAAAAACCAGTGAGGCCATTTCCGTGTGTAGTGATCCGAACTCAGTTACTATTGATGGAAATGAGGACTGGGTCATGGGGCGCAATGGAGTGAAGTAATATATACTTTAGCATACGTGTGCGTACGCCATATCAATATGCTAGTGAGGTGGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGGGTGTGTGGGTGTGTGGGTGTGGTGTGTGTGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGTGTGGTGTGGGTGTGGTGTGTGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGTGTGGTGTGTGTGGGTGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGTGT tpg|BK006940.2|:268423-270160 7X501=45S 24S3=362S 
 tpg|BK006940.2| 76774 + tpg|BK006940.2| 77153 - INS GTTAGCGTGTGCTACTTCAACCGAAGAAGAAGAGGCTTTTCAAGAATGCAAACGTGAGGTTGGCGCGCCCTCCTACAATTATTTGTGGCGACTGGGCAGCGACACTGAACATAGCTCTTGAACAAGACCCTTTTTTGGCTGCAAGGAGCAAGACTGGCTGGGGTTCCACCTCAAAGAGCCACGCTCTGCTTTTTTTCTATCTGTTTGTGTCATATCTATCTGTCTATTTATCTATATATATATTTTTTTAT tpg|BK006940.2|:76258-77669 7X2=325S 126=7X 
 tpg|BK006941.2| 529060 + tpg|BK006941.2| 529215 - INS CTTGGGGTCTTGATATAAGTACTCTTCCACTTTTAACTTACTCCCAGTTAGTATAATATAAGTAGTTAAGGTATGGCAAGCTGCAATCCGACCAGGAAGAAGAGCTCTGCTTCAAGCCTATCTATGTGGAGAACGATTCTCATGGCGTTAACAACACTACCGCTAAGTGTTCTTTCGCAGGAGTTGGTTCCAGCTAATAGCACAACATCGAGCACAGCTCCTTCCATCACTTCGCTTTCCGCAGTTGAGTCA tpg|BK006941.2|:528542-529733 7X322= 9S228=7X 
 tpg|BK006941.2| 988508 + tpg|BK006941.2| 988471 - INS TGAACACTATAGCATAGTCCAGCCTCAGCAGCCGCAACAAGTACTTTCTCCACAAGCATTATCTGGACCTCCGATGAAGAAATCAGGAACACTATCTTCGACAGATGATCTGAAAACAACTTCCTTGCCAATTGTTAATTACCCAATGCCGTATCATCCTGGAGCTTTTGCCCAGCAGCAGCAGCAGCAGCAGCAACCGCTCCCTACAGTCC tpg|BK006941.2|:988033-988946 7X302= 199=7X 
 tpg|BK006941.2| 15614 + tpg|BK006941.2| 15803 - INS TGGTGTTTGTAACGCTGTCTTGTTGCCTCATGTTCAAGAGGCCAACATGCAATGTCCAAAGGCCAAGAAGAGATTAGGTGAAATTGCTTTGCATTTCGGTGCTTCTCAAGAAGATCCAGAAGAAACCATCAAGGCTTTGCACGTTTTAAACAGAAC tpg|BK006941.2|:15288-16129 7X136= 123S3=56S 
 tpg|BK006940.2| 197698 + tpg|BK006940.2| 197045 - INS CATAAATCATAAATCCTCACCCTCTTTAAAGGGGTCCTCCTCACCCTCTTCATGTACTTTAGATAAGGGCAACTACGATTTTCCCTTTAGTGCTATTTTGCCTGGTTCGTTACCAGAGAGCGTAGAATCTTTGCCAAATTGCTTCGTGACATATAGCATGGAATCCGTTATTGAACGCAGCAAAAATTATAGTGATTTGATCTGTAGGAAAAATATTAGAGTTCTGAGAACCATTTCACCCGCAGCAGTGGAGTTATCAGAAACTGTTTGTGTAGATAACTCATGGCCCGACAAAGTGGATTATTCTATTTCAGTACCCAACAAAGCCGTAGCTATTGGTTCAGCCACCCCTATAAATATTTCCATTGTACCTCTTTCGAAAGGTTTGAAATTGGGCTCAATCAAAGTCGTATTA tpg|BK006940.2|:196201-198542 7X5=207S 10S393=7X 
 tpg|BK006941.2| 650103 + tpg|BK006941.2| 649949 - INS CCTTTGGTTGTAGATGGTGGTGGCGGTGGGTTCTGTAATTGAGAGGCGGTAGGTGCCCTGGAATTTCTTAAAGAGTAAGTTCTGTGCATACGATATACTTGATGCTGATATATTCTTCACTTTGCAATACTGCTAACAATGGAAAAGTATAGGTA tpg|BK006941.2|:649625-650427 7X4=73S 74S4=7X 
 tpg|BK006940.2| 83002 + tpg|BK006940.2| 83443 - INS TTGCTACAGATGTCTCAAGCAGTGCTAAAAGCAGTCTCAGAAGTAGATTATATGACCTATATCCTAGAAGGAAGGAAACAACATCGGATAAACATTCGGAAAGAACTTTTGTTTCTGAGACTGCAGATGATATAGAGAAAAATCAGTTTTATCAGTTGCCCACACCTACGAGTTCAAAAAATACTAGGATAGGACCGTTTGCTGATGCAAGTTACAAAGAGGGAGAAG tpg|BK006940.2|:82532-83913 7X179= 8S206=7X 
 tpg|BK006938.2| 866567 + tpg|BK006938.2| 866268 - INS TGCGGGAACGGATGCCCGAGCCCGTGCCCGCGCCCGAGCCTGCTGCGGTGGTACCGGGGGAAGAAACCGCTGGAGCTTGTGGTGGCGGCAAATGTATTTTTTTTTTGGCGCCGGCGACGATAGTAGTAGTGGCAGTGTTACTATTAGTGGAGGTGGAGGAGTAAGGGAAAACATCCTCGTTGGTTGCAGTATACTG tpg|BK006938.2|:865862-866973 7X98= 238S3=7X 
 tpg|BK006938.2| 63437 + tpg|BK006938.2| 63964 - INS TTGAAGATATCCACAAGTGAGTTGTTCAAATCACATTCTGAAATAAGTTCTGATGACGAATGCTTGCTGCTATTTGTCGATTTTGTAGATATGGTGCTTATCACACTTACCAAATCCAACGGTTTTATGTCCTCTAAGAATAGAGTATAGTTCCCGTGTTTTGATACATATAAAGCTTTACAACTTGAAAAACATAACCTTTCAAGGTGAATATCTCTCAGTATTACTGTTGGGGATGCGCCTGAGTCAGAATCTAAATCTGGCAGTTCAATAT tpg|BK006938.2|:62875-64526 7X71=66S 2S1=241S 
 tpg|BK006941.2| 50918 + tpg|BK006941.2| 51032 - INS ACATTCAAGTGGGTATGGGTATCTTCCATAAGTATTTGTCATATTCTAATCCTTTATTGGAAGACCCTGACGAAACTGAACATGCGTCTGTCCTAATAAAAGTAAAGTCCTCTATCCAGGAGCTGGTTCAATTGTACACAACAAGATATGAAGATGTCTTTGGACCTATGATCAATGAATTCATACAAATAACTTGGAATCTTCTGACCTCAATTTCAAACCAACCTAAATACGACATCTTAGTATCCAAGTCCTTGTCATTTTTGACTGCCGTAACACGTATTCCAAAATACTTTGAAATATTCAACAACGAATCTGCCATGAATAATATCACAG tpg|BK006941.2|:50232-51718 7X4=164S 103=1X64=7X 
 tpg|BK006941.2| 85626 + tpg|BK006941.2| 85900 - INS TGAGTAGACACGTTGGATCTTATTTGAAAATGATTACGGAACAAAAGCGACAAATCGAAGAGTTACGCGAACGTGAAGAGAAGATGATTTCTTTGAAGCTAACGAAATACAAACTAAACAAAGAAAAGATCCAGTTAGCCATTAACGAGTGCGTCAATCGTGTTCAGCAAACGTATGCAGGAGTGGAAACGTATCAAGTAGCCAAGACCTTGAAATCATTAATAC tpg|BK006941.2|:85162-86364 7X135=33S 6S1=156S 
 tpg|BK006940.2| 42023 + tpg|BK006940.2| 42665 - INS CAAGAAAGTGAGCGTAATAGGTAAAGTAAGGTAGAACGGAATAAAATGCTCAAGCGTATTGTTGGATTGCCTGCAAGGCGTTGCTTTCATAGAACGTCCTTTTTGCTGGGCAGTGACTTTGAAACTGTGCATATTCCCAATACGAACCACTTTAAAGATTTACTTATAGAGAACGGTAAATTTCAAGAGGATCAAGCAACTACAATAGTAGAGATAATGACAGATGCAATTAGGGGCGGGGTTAATCATGTTTCACAGGATCTGGCAAAGAGAGAAAAATTGACCCAACTTAGCTATCAACAACGTGTTGATTTTGCAAAGTTAAGAGATCAGCTATTGAG tpg|BK006940.2|:41327-43361 48S161= 171=7X 
 tpg|BK006941.2| 240243 + tpg|BK006941.2| 240449 - INS AATTTATTAAAATTGCCAGATTATAGAAACAAAACAATTTTGAGAGAGAAATTATTATATGCAATAAACTCAGGCGCCAGGTTTGACTTATCATAATTCCCAGAAGATTAGGGAGGTAATTAATTAATAGGCAGATTTCTAGTTCTTATATATTACTATAGATAAGGAAATTATACGCTTGTATGCAGAGATAATTTAAGTTTTGCTTTGTTCGCCACCATTCTAGTTATGACC tpg|BK006941.2|:239761-240931 7X5=112S 111S6=7X 
 tpg|BK006938.2| 38794 + tpg|BK006938.2| 38785 - INS GAACAAGGCCTTCTGTTGGTATATTTTCTTGAATAGGTTCTTCTCCATAGAATTGCCTCCTGAATTTAAATTCGAATGTGATTGGTCCTTCATTTCACTAAATTTCTTGATGAAGTGGTAAAGTTTTTTACGTGACATAATTGGATTTGGCAAGTATCGCGGTATCTTGTTTTTTGATCTGAAACAATTGGATAAAATGTAAAAAACGAAAATCACTGATGAGACACTATCTCTTCGTAGCGATAGTAAGGCTCTCGTGGTTTCAATATCAAAATCCTGATCCCAAATTTCAAAAAATGCACCTGAAATTCTCGCTTCAATGATCTTAGATAACAAAAATTGGCATGAATTGATTAGACTTGCGTACTTCTCAGGATTGAAGTTGGAAATAATGATTGGCTCATGACGGGCTTTCTTCAAAAGTTCCCTGATTG tpg|BK006938.2|:37903-39676 7X186= 217=7X 
 tpg|BK006940.2| 220371 + tpg|BK006940.2| 220723 - INS TGTAACCGACCAGCCTTCAACAATGGTTTGTCAACTCTACCACCACCGGCAATGACACCGATGACACCTCTGGCATCAGAAGAGATAACCTTCTTGGCACCGGATGGTAATCTGACTCTAGTCTTGTTTTCGTCTGGGTTGTGACCGATGATAATAACGTAGTTACCGGAAGCTCTGGCTAGGGCACCTCTGTCACCTGGCTTTTCTTCAACGTTGGAGACAATGGTACCTTCTGGGACAGAACCCAATGGCAAGACGTTACCGACGTTCAAAGAAGCCTTCTTACCGGCGTAAATGAATTGACCAGTGTGGACA tpg|BK006940.2|:219727-221367 7X186= 158=7X 
 tpg|BK006940.2| 60175 + tpg|BK006940.2| 60239 - INS TAGGGCCAGAATTTAGATCCGAGCAGGTGTTGAAAAGCGAATCTCAAGCGTTCAGAGATGTTAACAAGAAATCACCAGAATTCAAAAAACTGGTACAAAATGCTAAATCTGTATTCAGATCATCTCAAATTGAGCAGTCGAAAATTTTGTGGCCTCAGAGTATTAGGGCCAGAATCGGTTCGGTATTAATCTCAATGTTGATTCAAGTCGCTAAGGTATCTGTGCAAGGTGTTGACCCTGTGACAAAAGCTAAGGTTCACGGTGAAGCTCCAGCTTTTGCGCATGGTTATCAGTACCACAATGGTTCCAAATTGGGTGT tpg|BK006940.2|:59523-60891 15S153= 9=1X290=7X 
 tpg|BK006940.2| 28910 + tpg|BK006940.2| 29387 - INS TTTTTACGACAAAGTGTCAGTGTGCGCTTATCACGCTTCCTCTTTCTAATCCGCTTGAATCGACAGATGGTTCTAAAGAAGATGTAGATGCGCTTCCTTAAGTAAACACATTGCTACTTGCATTTTACCTTTCAAGATGTAGTGATTACGGACAGTTGAAGAGGCTAATAGCATCTATTTCTTCTTTAGTATATGGTTCCTGCAGGGCAAACAATTATTTCCTTTGCAATTTTGCGGCAGTGGGGAAGAATGATAGCACTAATAGTG tpg|BK006940.2|:28362-29935 7X13=89S 134=7X 
 tpg|BK006941.2| 136126 + tpg|BK006941.2| 136490 - INS CTATGGTGATCATAATGGTGAATTCTCTGGTAAATTGGTCGATGTACTTGGCCAAGACCGTCGTGATAGAATTTTAGCCGCATTATTTGTATGCAGGAACGACACTTCTGGTATCGTACGTGCTACGACGGTTGACATTTGGAAGGCATTGGTTCCAAAT tpg|BK006941.2|:135792-136824 7X8=72S 71S9=7X 
 tpg|BK006941.2| 256366 + tpg|BK006941.2| 256795 - INS AATAAAGGAAAATTATAGAGGAAAAAAAGTGTAGAAATAGAAAAAAAATAAAAAGGATAATACCGATCAGAAAAATCCTCTTTCTTGCTCTTCTTCTTTTCTTTGTATTTCTCCTGAAAAAATTCAGAAAAACATATATTGGGTTAAATACATAAC tpg|BK006941.2|:256040-257121 7X6=72S 73S5=7X 
 tpg|BK006940.2| 192109 + tpg|BK006940.2| 192884 - INS AATAAGAGTATTCTGAGAACGGTACTGATTTGATGACACCCGAAGATCTTCCTGATTTGCTATCAGATGGTATAGTATTATCTTTTGCTAATACTACAGAAACGGGCTCGGATTCGGACTCCACGTTAATTGACAGTGAAGATCTTCGGAGATGTATAGATATGCCGGACCGCTCATGCTCTGCTCAACGAGGCAATTTGTGTTCATACAGTTTTTGGGATATTCCTTTCAGTTTCTTGAATACAGTCCATGATATATTCGGCATGACTAATATGGGTAATTGCGCAGTTATGGCT tpg|BK006940.2|:191503-193490 7X6=258S 148=7X 
 tpg|BK006941.2| 483059 + tpg|BK006941.2| 483237 - INS CAAAGCTGAGTTAATCTCGGAAAATCTCTGTGTCCTTCCTTTTTCTTCTAGCTTCCGTTCCGAGTCTCATCTTCTTTCCCGTGCCGTCGGGTTTAGTAAAGAAATGTAAAGAAAAAATGTCGTATCGTACCCGAGAAATATTTCAATTCTCTTACGTATGCGATAGCAGTTGGAAAGATCTGATTCGTTACGATGACTTGATAAGCGCGGGCTTTTTCGCCCTATACGGCTT tpg|BK006941.2|:482581-483715 7X59=57S 1S1=403S 
 tpg|BK006941.2| 475334 + tpg|BK006941.2| 475641 - INS GTTCACTACCATACCAATTGTTCTTGAAATACAAAAAATATACGAAACAGTAGTTGGATCCAACAGTTTATCAGGGACCTTTTTCTGACTTATCACCACTGTACAATCTTTACCTCTGACCGCTAGTGAGTTTATGTTAGTTTGATTAGTCGCTTTAAAGG tpg|BK006941.2|:474998-475977 7X4=199S 81=7X 
 tpg|BK006941.2| 87477 + tpg|BK006941.2| 87553 - INS CCCCCTCCCCCCAACAAACCCCCCTTCATATAGAAATGGCTAATACTTTCAAGTATTATCCTGAAACGATGGGTAATTCTAGTGGTTATCCAATTAGTTTGCCTTTTCCGAAAGGTTCGGCTACTTCTGCTGTTAATGTTGCTAGGCAACTGCCTAAATATTTAGGTCATGTTCCCTCGCAATCAGTTCATACTCAGTTGCCATCCATGGCTTCTTTAGGTTACTTCAATCAGCCAAGTTCTACTTACTATGCTCCTCCTGCACCACTTCAACAGCACCAGCAACCACCTATCCTTCCCCCTCCGGGCCTAATGTACAC tpg|BK006941.2|:86825-88205 7X260=19S 2S1=268S 
 tpg|BK006938.2| 1407380 + tpg|BK006938.2| 1407642 - INS TACAATACAGTGTAGGGTTACAGTTCGAATCATTAGATTTTACTTTTCTGAGCGAAGATGAGCTACTGACTTTCCTCAAAGATGAATCCTTATTACCAGAACTCACACTATATGACTTTGAAGGTGCCAAATGGGGAAGGCCTGGAACGGACAACTGATCTGTGTCACGATGATGGTGATGATGATGTTGTTGTTGCTGGTCCCCTGGGCTGTCTAGCGAGTGCCTAGATTTAATAGCACCCAGTGCAGCATTGCCATCTACATTCTTGACACTCGACGCGAACTTGATTTGCGGAGAACGTGATCTCGACGCACTCGCACTTGAGTTTATATCGGTAGCAGTAGG tpg|BK006938.2|:1406674-1408348 7X310= 232=1X92=7X 
 tpg|BK006938.2| 1222061 + tpg|BK006938.2| 1222506 - INS AGAACCTTTCGGAAGATTTTGTTAAGATATACAAACAGTTTTTTCCATTTGGTTCTCCTGAAGATTTTGCTAATCACCTTTTTACAGTTTTTGATAAAGACAACAATGGATTCATACATTTTGAAGAGTTTATCACAGTTTTGAGTACAACGTCCAGAGGAACTTTGGAGGAAAAACTGAGCTGGGCTTTCGAACTTTATGATTTGAACCATGATGGATATATTACATTTGATGAAATGCTAACCATTGTGGCGAGTGTTTATAAAATGATGGGGTCTATGGT tpg|BK006938.2|:1221481-1223086 17S131= 63=86S 
 tpg|BK006938.2| 234743 + tpg|BK006938.2| 234610 - INS GGTAGCTATAGAATCTAGCATCGACCACAGCTTCCATTATCAAAATTAAGAAGACGAATAGTATGATAGATATTGCATTGCCAGCACCACCGTTGACTAAATTCATCAACAGACTGATCAAGCATTCTAACGTTCAAACTCCGACTCTGATGGCTACCTCTGTATATTTGGCCAAATTAAGATCAATAATACCGAGTAACGTTTATGGTATAGAGACCACCAGGCATAGAATATTCTTAGGTTGCCTAATATTAGCTGCAAAAACGTTAAATGATTCCTCCCCTCTTAACAAACACTGGGC tpg|BK006938.2|:233994-235359 7X215= 283=7X 
 tpg|BK006940.2| 175439 + tpg|BK006940.2| 175573 - INS CGCTTGGTCTGTTTCAATCAAGTCTTCCATGTAGGCACCGAACCCAGAAACGTTTGTTGTGATAGATGGGACACCCATGACGGTACATTCTGCTGGCGTGTACCCCCATGGTTCGTAATAGGATGGAAAAACACCCAAGTGACAGCCGCGAACAAACTCGTCATAATCCAAACCAAGGATAGGGTTATTGGCGTTTAAGAATTCAGGATGGAAAATCAATTTT tpg|BK006940.2|:174979-176033 7X5=106S 106S6=7X 
 tpg|BK006941.2| 951286 + tpg|BK006941.2| 950588 - INS TCCCAAATGTTCACTGGTCCAAAAATCGATGTGTCTCCAAGCTAAGAGGGTTTCAGAGACACCATCGTTTGACTCCGTGGACGTAAATTCATCAATATTTATGTCTTCATTAGATGGCACGCCATTTTGAAATCCCATGCTCATTTCCTCATCTACACTATTCAAATGCATTTGAGAGGGATTTACCTGACCATTGTTGCTGTTTAAACGTTTACCCATGTTAAAAGTAGGCGTTTCATCGGGGTTATACTCTGCATAATGGTCGTCAGTGCTGAGGGAGTATACCCATTC tpg|BK006941.2|:949992-951882 7X5=300S 146=7X 
 tpg|BK006940.2| 258876 + tpg|BK006940.2| 259216 - INS GAATGGAAGCCACAGCCAACAGGCACCTACATGTTCGTTATCCATTTTTGAGGAAAAAATAGAAGTGATAATAATAATTTTGCTCGAACTACTCGTAAAGCTACTTGAAAAACGGCTCGAGATTACGGAAGAGTCGGTAGTAAACCGACTCTCAGTGTCACGGAATGGAAGCGCCTTGAAACTACTAATATCAGGTATGCATTGAGGGGCAAGGCAACCTGAATATGCAAAGAGCATAGTCTTAACTTTCGTAGTACGTAATACTTCGGCATTAATTTGGCCTACCGCTTTGCCACAGTTGAGTGGTCACTGGAGTATTAGC tpg|BK006940.2|:258218-259874 7X5=183S 302=7X 
 tpg|BK006938.2| 104740 + tpg|BK006938.2| 105321 - INS GGGTAGTTCGGGTAGTTCGGTTGGCGAGTGGACACGATTTTTCGCTACCAAGTTTTTGGAATATGCCCAAATGGTGTTTGCGCTGGGCTGGTGGTAGCCGTTGAATTAATGATTGCACGTAACTCTGCAGTAGCTTGATGGTATTATTTTTTCTTTCTAAATGCAAGTGGGTAGTTCGGCTCCTCTCATCGGCCATTTTCTTATGCAACCTTAGATCTTGCAATTCCTGTTCCTGGATAGCGAACAAATCCTCTGGATTGTTTTCCTCAAAGGGGTCCACCAAAGTCACATTGGTGGGGATTTGTACTTGATTTTGTGTTTCTGTTTCTATTTGCCCCTTTGTTTCTGATTGTTGCGATAGTTCTGCTTGTAATGCTTCGATAGTCTCCCTCTGGTTAGCGATGCTTTTCTTGTAGGATAACATCGTGAGATTGGCTTTGTCGACCAGCTCAGGAA tpg|BK006938.2|:103814-106247 7X199= 8S434=7X 
 tpg|BK006938.2| 900359 + tpg|BK006938.2| 900559 - INS ACCAACGACTCAATTACCTAGAATCCTTTTTAACAATTTCCTTCTTTTCGGAGCTCGATTCTATTTCGTTATTGTACACTTCAGTATGCGTATTTATGTCCTTTTCGTCATCAGTATGTTTCTTCGGAGACAGAACATTGGTCATTGATTTCCTTCCCCTAATGGGATGTCTCAAGTACCTATACGCGTCGCCTTTATTTTTCTCATTATCTTCTAATATGATCTTCGCTCTTTTAGCCCACTCGCTTAGGTCAAGAC tpg|BK006938.2|:899829-901089 7X259=1X167= 1S241=7X 
 tpg|BK006941.2| 974007 + tpg|BK006941.2| 974594 - INS CCGCTATCAAGAGTAGTACGGCCTGTTGAGAACAAAAAACTGTAGTATCTATCGCTCACTATATATCTATTAAGTTAGGATTTTCTTGCTGATGCTGCTGTTGTTGCTGTTGTTGATTGATGGGGACAAACGCAGTGGGAACCATAACATACCCTGTTTGCTGACCCTGCATCATTTGTGGTTGCTGCTGCGCACCAGTAGAG tpg|BK006941.2|:973587-975014 7X8=4S 5S181=12S 
 tpg|BK006940.2| 198392 + tpg|BK006940.2| 197828 - INS GTGTAGATTGTGAGATTGATACCATCCTGCAAATCCCGAACAGCTTATCAAACTGTGTGCAAGATTGTGATGTCCGCTCTAACATTAAGGTTCGCCATAAGCTCAAATTTTTCATCATCCTAATTAACCCAGATGGTCATAAATCTGAGTTAAGAGCGTCCTTACCGATTCAACGTTTTATTTCACCATTTGTGGCACTTTCAATAAAACCATTGTCATCCTCGAATTTGTATTCGCTTTTTAGCACCACTAACCAGAAAGACGAAAACTCATCACAAGAAGAGGAAGAGGAATATCTGTTTTCTAGATCAGCATCAGTCACAGGGTTGGAATTATTAGCGGATATGCGTAGCGGTGGCTCTGTTCCTACCATTTCAGACTTGATGACGCCCCCAAATTATGAAATGCACGTATATGATCGTCTTTATAGCGGTTCTTTCACTCGCACGGCTGTGGAAACGTCTGGAACATGTACTCCTTTGGGAAGCGAATGTTCGACTGTCGAGGATCAGCAACAGGATTTAGAAGATTTACGTATACGGTTGACAAAAATTAGAAATCAACGTGACAATCTAGGGCTACCACCGTCTGCCTCGTCTGCTGCCGCTTCCAGATCGCTATCTCCATTACTAAACGTTCCAGCACCAGAGGATGGCACGGAGAGAATCTTACCTCAGAGTGCTCTTGGTCCCAATAGTGGCTCTGTGCCAGGAGTACATAGTAACGTATCACCTGTTTTACTT tpg|BK006940.2|:196328-199892 7X5=248S 163=1X568=7X 
 tpg|BK006941.2| 317296 + tpg|BK006941.2| 317427 - INS CAGTATATATAGCGAAGCTGTTATGGAGTTGAGAAAGAGATTGTTGGGGAAGGGACAGAATAAGGGTTTAGGATATGAAACTACGAAATCAGTCGATAGGCAAATTGAGGACCAGGACACGTTGCAACAGGATTTGATTCAGGATATGAGCAAACTTGTGGGCAGTTTGAAGCAAGGAGCTGTGGCATTTCAATCAGCACTTGATGAAGATAAGCAAGTTCTTGGA tpg|BK006941.2|:316830-317893 15S105= 101=19S 
 tpg|BK006938.2| 302861 + tpg|BK006938.2| 303583 - INS CGTATAGATGAAGTCTTCTTGGTGTCGCCAAGAAGCTTCTTTTTGTTCACACCGTTATTACCCTCAACGCCTGTGGGTACGATAGAGATGAACTCTATTGTCGAACCGGTTAGATCGATCGCTAGAAGAACGCCTGGAGAAGTTCACTACATTGAGGCGGAAGCGTTGGACGTTGATCCAAAGGCCAAAAAAGTAATGGTGCAATCGGTGTCAGAGGACGAATATTTCGTTTCGAGCTTAAGTTACGATTATCTTGTTGTTAGTGTAGGCGCTAAAACCACTACTTTTAACATTCCCGGGGTCTATGGCAATGCTAACTTCTTGAAAGAGATTGAAGATGCTCAAAATATTCGTATGAAGTTAATGAAAACCATAGAACAGGCAAGTTCATTTCCTGTGAACGATCCGGAAAGGAAGCGATTATTAACGTTCGTGGTTGTTGGAGGGGGCCCTACGGGGGTTGAATTTGCCGCCGAACTGCAAGATTACATCAATCAAGATTTGAGGAAGTGGATGCCCGACTTAAGTAAAGAAATGAAGGTTATCTTAATT tpg|BK006938.2|:301743-304701 7X274= 2S73=1X459=7X 
 tpg|BK006940.2| 75672 + tpg|BK006940.2| 75487 - INS CACACCTTCACCTTGACGAGTACAGGGATTTCCAGAGCACGAGGGGCGCTTCACTGGACACCAGGGCCAGTTCGCACTCGTCGTCTGATACGTTCACACCTTCACCTCTGAACTGTACAATGGAGCCTGCGACTTTGTCGCCCAAGAGTATGCGCGATTCCGCGT tpg|BK006940.2|:75143-76016 7X2=170S 145=7X 
 tpg|BK006941.2| 1036676 + tpg|BK006941.2| 1036802 - INS GTTATATTGCCTGTAAGAGGTGGTGAAATTATCATGAATGAAGAAATGTCGCAGCAATCGAGGTACTCCGTTGAAAGCACTTTTACCGATGAATTCGAATTACCGATGTGGGATCCACATGTAAAAACATTTTTATTACTTCAAGCTCATTTAAGCCGTGTAGATTTACCGATTGCAGATTATATCCAGGATACCGTATCAGTTTTGGATCAATCTCTACGTATTCTACAGGCTTATATTGATGTCGCCAGTGAATTGGGTTACTTTCATACGGTATTGACCATGATAAAGATGATGCAATGCATAAAGCAAGGGTATTGGTATGAAGACGATCCTGTTAGTGTACTTCCAGGATTACAACTGAGAAGAATCAAAGATTACACTTTTAGCGAGCAGGGGTTCATTGAAATGACGCCGCAGCAAAAGAAGAAAAAGCTGTTAACC tpg|BK006941.2|:1035774-1037704 7X220= 222=7X 
 tpg|BK006940.2| 184667 + tpg|BK006940.2| 185308 - INS GTTACTGCTATCCAATCCCAGCAACAAAGCAAGGCGGATCGCTGGAAATCTCATTCGATTCGGAAAACGATAGGGCTTTGCATTATCAAGATGACAACCCCGGTCGCCATCATCACCTCGATTCCGTGCCCACAAGGTACACTATCAGAGATATGGACAATATATCACATTACGATACCAACTCTAATTCCACTTTGAGGCCACATTATAACACCAATAACAGCACTATTACCATCAACAACCTCAACAACACTACTTCCAACAACAGCAACTATAACAATACCAATAGCAACAGCAACATCAATAATCCTGCGCATTCCTTAAGAAGGTCTATTTTCCATTATGTAAGCAG tpg|BK006940.2|:183949-186026 21S162= 163=20S 
 tpg|BK006941.2| 559979 + tpg|BK006941.2| 560028 - INS AAGGCTTCGTCACCTTCCGAGAGAATAGTCGAAATATGTTTAGTCCCTACACAAATTGCTAGACTACCTGTTTCGAGTTTCCTCTATTCCTTTGCTAACGGAGCTGCGGTATATAAACCATCGTAGACTCAAAGCCGTTACCCGACAACTATCGGGTATAGTGAAATGCCTATGTTTTCACTTTAAGACCTTAGAAAACTATCATGAGATCTCGCCTTCAGATGCAGATATTTCA tpg|BK006941.2|:559495-560512 7X1=1X8=4S 5S211=12S 
 tpg|BK006938.2| 358103 + tpg|BK006938.2| 358480 - INS GCAGATCTGCAATTGGAGGAGCGGATAAAGCAAGTTTCCCCCCTCAATGTAAATCATCTTAAGCAAAATTTTAAAATCTAGGCACATATAAAGAGAAAATGGGAATGATTTTGCTGGATAGGCTACAGTGTTAGGAATGCAGAATTAGGAACTATAGATGATGCGATTAAAGATATTAAACGAGAAGTGACAGTGGTGGCTTCGACAACGGCAGTCGTGCTCGGTCGACAACGTGTATGTTTTTGCCGAGCAGAGCAGGGAAAGTCCTTCTTTCTGCGCGTGAATCAAAACACATTGGTATCGAATTTAACATATCTGGGTGAGGAATGGACAATCCTAATAAAGTACTGGAGGTTTGTCTGTATTTCCAAGTTCTTGCTTGTAGAAACTGCTTTCTTTTCTCTTTTCCTGCAGCGGTCGAACATATGTGATTATTGATTAGCCATTTGTTCCAAGTCATATAGTAGTATTACGTGTTCAGATGCGGTGTTAGCGTATCTTTTTGTTAAATAAAATATCATTGTGCCGTTGCCGCCCTACCTGCCAAGGGTCAAAGAAGGCACCTTTATACGATGCCACCTTTTTATAGTATTCTACTACAGAGT tpg|BK006938.2|:356879-359704 7X335= 587=7X 
 tpg|BK006940.2| 199114 + tpg|BK006940.2| 199417 - INS GGAGTACATAGTAACGTATCACCTGTTTTACTTTCAAGATCCCCAGCCCCAAGCGTGTCAGCCCATGAAGTGTTACCAGTGCCCTCGGGCTTAAATTATCCAGAGACTCAAAACCTGAACAAGGTTCCATCGTATGGCAAGGCAATGAAATATGATATCATTGGTGAGGACCTTCCTCCTTCCTACC tpg|BK006940.2|:198726-199805 7X5=88S 90S4=7X 
 tpg|BK006941.2| 210544 + tpg|BK006941.2| 210688 - INS GAAAAAAACTCTTGCAAGTTTGACAATTCTAAGACAAAAAAACTACTGGGATTCCAGTTTTACAATTTAAAGGATTGCATAGTTGACACCGCGGCGCAAATGTTAGAAGTTCAAAATGAAGCCTAAGTATCACGCTAATTGAAGTTTTTTTT tpg|BK006941.2|:210226-211006 7X5=71S 71S5=7X 
 tpg|BK006940.2| 202061 + tpg|BK006940.2| 202135 - INS GTGTTAGGTCTTGTGTTAGGTCTAGTGGAGGAGGCATCTGTAGAACTGAATGAACTAGGAATGTCATTATAGTAATCGTCGTCGTCATAGTAATCGTCTTCGTCGTCATCGAAACTGCCACGACCACCGTTGGAGGGTCTGTAATTAAACGCCCTGGACTCTAAAACACGAAACAATGGATCAACTGCTGGAGGCGGTCTTATCCTACCAGACAAAATCATTTTCGCGGTACAATTGTCACCATAAAATTTTCTGTTAGCCTCTCTTCTTTCTATAATAGCCGAACCTTCCACAGAAACC tpg|BK006940.2|:201447-202749 15S24=1X117= 54=103S 
 tpg|BK006941.2| 944936 + tpg|BK006941.2| 945470 - INS GCTTATAAGTACCTTTGACTTTAGTACACTCTCGCCCGATGTTGCCCGTTATTATATCGCTAATTCTAACGCAAGATCAGCTTCCCCACAAAGACAAATCCAAAGACCTGCTAAACGAGTAAAGTCACATATTCCATACCGTGTATTGGATGCACCTTGCCTGAG tpg|BK006941.2|:944592-945814 7X10=10S 138=14S 
 tpg|BK006938.2| 200662 + tpg|BK006938.2| 199941 - INS GGTTGTAATTGGAGGTGCGGCAAGTGTGCAAGACGGGTAAAGGAGAGTATAGAACGATGTCTGCTAAAGTTCCATCTAACGCCACGTTTAAGAACAAGGAAAAACCTCAAGAGGTTCGCAAAGCCAACATCATCGCTGCACGTTCTGTTGCAGATGCCATCCGTACTTCATTGGGTCCCAAGGGTATGGACAAGATGATTAAGACATCTCGTGGAGAAATCATCATCTCTAATGATGGCCACACCATTCTAAAACAGATGGCCATTCTGCATCCGGTGGCCAGAATGCTAGTAGAGGTTTCTGCCGCGCAGGACTCGGAAGCCGGTGATGGTACCACTTCTGTGGTGATCTTGACCGGAGCTCTATTGGGTGCTGCTGAGAGGCTGTTAAACAAGGGCATCCATCCAACCATCATTGCGGACTCCTTTCAAAGTGCTGCGAAGAGATCTGTCGATATTCTTTTAGAAATGTGCCATAAGGTTTCGTTGAGCGATAGAGAAC tpg|BK006938.2|:198925-201678 7X5=371S 251=7X 
 tpg|BK006941.2| 505516 + tpg|BK006941.2| 505994 - INS TTTTACGTATAGAATCGACCTTTGGAAAGGGCCCCAATGGAAAGAACTTCAATGTTTTTTCCTCTACAAGTAATAAGAGCATAAAATGGACCTAGATCTAGCCAGTATCTTAAAAGGTGAAATTTCTAAGAAGAAGAAAGAGCTGGCCAACTCTAAAGGTGTTCAGCCACCATGCACTGAGAAATTCCAGCCACATGAATCCGCAAACATAGACGAAACACCGCGACAGGTAGAACAAGAAAGTACAGATGAAGAAAACCTGTCAGACAATCAGAGTGACGATATTAGGACCACCATTAGCAAATTAGAAAATCGGCCAGAAAGGATACAAGAAGCGATAGCTCAAGACAAAACCATC tpg|BK006941.2|:504786-506724 7X264= 336=7X 
 tpg|BK006938.2| 851377 + tpg|BK006938.2| 851564 - INS TTCATGGTTTCCAGGATTTGTTCTTCACTGAACTGGAGAAATTGATATTGGAGAGTTGTACCGAGCCATTATTGGCAGTATATGATTGCGTATATAAAAAGGAACTTTTGAAAATCCCCGGAGCACAAGATATAATAAAAAAGTTGATTAGTGAGCAGCTGTCAATTATCGATCGATCCTACCCGTCACTAAACACCAACCC tpg|BK006938.2|:850959-851982 7X49=52S 1S1=160S 
 tpg|BK006940.2| 70704 + tpg|BK006940.2| 70868 - INS CGATATCGTCTAAAAGTAATTCGAAAAATATACAACCAACTGACCACCAGTCGCATTGCTTGTTATCTTCACCCTTTCCTTCAATAGTTTCTGGAGCGAGATAATCGGGAGTCCCAAAAAATTTCTTATTTTGCTTGCTATCATCAGGATAAAACAAAGCTAAATCCGAAGGTGCTGGCGAAAGGGAAATGTTATTATTCGAGTTAATATTCGTATTGGTAGCTGCGATAGCATCTGAAGATAATAGGTCATTAGAAAAGGATTTATTC tpg|BK006940.2|:70152-71420 7X203=1X154= 253=7X 
 tpg|BK006941.2| 582398 + tpg|BK006941.2| 582568 - INS GTACGTGGTATGGTACTGACTTTGAGGGTACGTGAATCATCGAAGGAAACATAATTGCACTGATATGTAAACTTCCTAGTTTCAAATGTGTTCTCGGAATACCAAATAACCTCTAGCCATAAGTTTATTTTCAAACTTTTTCCTCTTAGGTGATAAGGGAGATTAGAAAAAAAGAAATATTTATTATTGAAATAACTGTCCAAAGAAGCAAAGTGAATATAGAAGAAAAAATGCGAGTACTTACGATTTTTTATTTAGCTAAGTAACCAACGTGGTGCCATATTCACGACATAGCAAGTGTCCATAGTTGCATGCGTTTTCTTTAATATCATTGTGTTTTATTTTTATTACTTTAAGAAAAAATACAGTAGCTTTCATGCCTGCACAAATTTAACAAGAGTTTCATGGGGTACATTTTTAATGCCTCAACTATTTGGTATTGTTC tpg|BK006941.2|:581494-583472 7X288= 76=1X355=7X 
 tpg|BK006940.2| 157495 + tpg|BK006940.2| 157598 - INS TAATTGATGCAGGTGCAGAATGGAGACAATATACAAGTGATATCACCAGATGTTTCCCAACTTCAGGCAAGTTTACTGCGGAACATCGTGAAGTTTACGAAACCGTTCTTGACATGCAAAACCAAGCAATGGAAAGGATTAAACCTGGTGCTAAATGGGACGATTTACATGCACTGACA tpg|BK006940.2|:157123-157970 7X4=18S 17S140=7X 
 tpg|BK006941.2| 575353 + tpg|BK006941.2| 576027 - INS GTGCAACAATTCATGCGGATGCATTTTGGCTGAAATGGTCTCCGGGAAGCCTTTGTTCCCAGGCAGAGACTATCATCATCAATTATGGCTAATTCTAGAAGTCTTGGGAACTCCATCTTTCGAAGACTTTAATCAGATCAAATCCAAGAGGGCTAAAGAGTATATAGCAAACTTACCTATGAGGCCACCCTTGCCATGGGAGACCGTCTGGTCAAAGACCGATCTGAATCCAGATATGATAGATTTACTAGACAAAATGCTTCAATTCAATCCTGACAAAAGAATAAGCGCAGCAGAAGCTTTAAGACACCCTTACCTGGCAATGTACCATGACCCAAGTGATGAGCCGGAATATCCTCCACTTAATTTGGATGATGAATTTTGGAAACTGGATAACAAGATAATGCGTCCGGAAGAGGAGGAAGAAGTGCCCATAGAAATGCTCAAAGACATGCTTTACGATGAACTAATGAAGACCATGGAAT tpg|BK006941.2|:574369-577011 7X10=16S 470=7X 
 tpg|BK006940.2| 136018 + tpg|BK006940.2| 136303 - INS GTATACTGTTCTTATCCAATTTATTTTCTACAAGTTCTAAACCTCTGACGGTTTTAGAATCAATCAGCATTGTATTTTCTGTTCCTTCAAACTGTATACGTAGTTTTCGAAACGCATTCAAATTTCGGCTGCTTTTGGATATAATCTCTTCCATGTAGCTTATCGCAGCAGATGCAGCACAAAGAGCAAACGTTTTATCTATAATCTCCTCGATTTTCAAGTCCTTTTTTGTATCATCCATTAAATACTTTGTAATCGCCGCCAGTCCATCTTGGCTATTGAAGCACTTTCGTGAACCCTCTTCAATTTTAACTGTCTCGGCCACATTAAATTTTATCATTGTCGCTAATTTTGATACTGTGGGAGCT tpg|BK006940.2|:135268-137053 7X6=46S 338=1X6=7X 
 tpg|BK006940.2| 236699 + tpg|BK006940.2| 236713 - INS ATTCTTAACACATCCTTGGAACAATTTTTGGCATAATGTTATATTCGACATAATTCAGCAAATCTTCAATGGAAGAATGGATTTTTCCTATAATTCCTTCCTTGTTTTGTCTCTGTTTAACTTAAAGAGCTCCTATCAATTTATGACTGATATCGTCATATCAGATGAAAAAGGAACGGATGTTTC tpg|BK006940.2|:236313-237099 7X3=246S 93=7X 
 tpg|BK006941.2| 631501 + tpg|BK006941.2| 632136 - INS TTATTAGACGAAAATCGGATTCACTAAGTGATTCATTTTCTAAATGAGAGTTGATAGACTTGAAGAAAGGAACTAAGTTTGCAAATTTTTCTAAGATACTCTTCAAAGCTGAAAATCTATCGCAGTTACAGGAAAGGATTGAAGTAAGTTCATTGCAGTTAGGTTGTGTATAATTTTGGCAGTATAATAGGAAATCCGATTTTAGGGAGTCGTTTAAG tpg|BK006941.2|:631051-632586 7X129=34S 8S1=188S 
 tpg|BK006940.2| 256118 + tpg|BK006940.2| 256610 - INS GAATAGTGGGGTTCAGGGGCATAAGAAGCTCACACAATGCGGAAAAACAAAAGGGGACTGCCATTCTTCCTGAAACCCACGCGTCACTGCTATACTGAGATCTGGCCAGGGGCAACCAGTATACTTAGTGGATAAACGACAGGAACACGTACTCCTTAAAAGCGTCTAAATCTTCATTTTTCCGGTTTATTTCCAACCGGGAAATAAATTATTCCTAATAAAATTTCCGGGGTTTGCAGGATGCGGGGTAAAAGTAAAAAAATGAAAAAGATGTAAAAAGAAA tpg|BK006940.2|:255538-257190 7X1=193S 266=7X 
 tpg|BK006941.2| 592069 + tpg|BK006941.2| 592064 - INS AGCTACTGGTGCCTTTGGACTCAGCTACTATCTAGCTGCACCAGGAGAAAGACCAAACTACCTTTTGTGCGGACTTGGTGTCGCCCCATTATCTGCAGCCTACCTATACTTAGTATCACTGTTCAATCACAAGCTAGCCCCAAAATGCACACGTGACCAAAATGATTTAGAAAAGCAAAAGGATGAAAA tpg|BK006941.2|:591672-592461 7X5=89S 89S6=7X 
 tpg|BK006938.2| 948339 + tpg|BK006938.2| 947782 - INS CTCCTAGTAGTTACGGCGTTATTGATCCTCCGCCCAGTGACATCAGGGCTTTAAAGACGTGCGAAGACCTAGTTAATAAAACTAAAGGAATGAAGGCAGTTAAATGGGAGCCTTCCAGTGAACTGAGCAGGGAATTGTTTGATCTCGCAAATGAAGCAGATGTTGCTGACTCAGGTAACGAGATAAAAAACGAATTCGAAATTTCCGGAGAACCACTCCTAGATATTTTAAAACCAATGGTTTTGGAAAACGGAAGGCCCCCATATACTGTTAATGAATGGTGGGATTTGACCAAAAGAGTTTATAATGCACAACAATTAATGAGAGATTATTACCTTTCTTTCCCGG tpg|BK006938.2|:947072-949049 7X5=342S 327=7X 
 tpg|BK006938.2| 956299 + tpg|BK006938.2| 956774 - INS GGATACAGAAGAATATGTCCTACCGCTTTCTTTCCAAGTCTGTTTATGAAAAGTTCGTTAGCCCCGTCGATAACACGAATGAGAATTTGTCTCCAAAATCCTACGTGTACATGCACGATAGTAAAGCTGCCAAGAATTTATCTTATACATCTTCAAGTGAGGAAGAAGATGGAATCAAAGAAGGGATAGACGATGATAATGGCAGTCGCAGTGGCAGTTTCGGAAAGCTAGACACAGACACTGGATTGCATTCTTCGTTCAC tpg|BK006938.2|:955761-957312 7X278=12S 12S197=1X36=7X 
 tpg|BK006940.2| 133575 + tpg|BK006940.2| 134326 - INS TGAAGAAAGCCACCTAATGTAAAACTCTGTACAGAAATAATGGATTATAGTTTTAAGCTAAGCGGAAAAGCCAAATTATTCTTCAAAATTTTCGATGAAGTCGGAGTTTATTTCTTTTAATTTCCCTAAAGTCAAGGGCTCTTTTTCATTTCCTGCACATTCTTTCAATATCGCTACAAGATTGTGTAT tpg|BK006940.2|:133183-134718 36S111=9S 166=7X 
 tpg|BK006941.2| 750111 + tpg|BK006941.2| 750055 - INS GAACGTAATACAGACATTTCCGTGTAGAATGACAAAAAAGCTAGAATATTACTATATTTTCCTTAAAAGAGCAATATTTGCGATGAGGGGCTCTCAATGACAATGTTTGACTTCTCTATTGAACTGTAAGCGAAGCAAAACCATATCTTGTCAAAGTATTCGAAGAATGGATTTTTACAAATTAGACGAGAAGCTGAAGGAGTTGAAAAGGAAAAGAGTAGATGTATCTATAAAGAGTAGGAAGTTGGCTGACAGAGAGATTCAGGAAGTAAGCGCAAATCGAAAACCAAGAGTATACAGTATGGAAGACGTAAATGATGCAGATGAATCAGTAG tpg|BK006941.2|:749371-750795 7X270= 168=7X 
 tpg|BK006940.2| 63322 + tpg|BK006940.2| 63994 - INS TGATATATGTATACATTCATCTTCAGGGGTGACTTGATAGAAAACCAATTTGTATTGGTTTTGCCTTATAGAGACGAATCTGATCCAGTCTCTTAGCTGATTCTTCTTCAAATACTTCTTTGTTAGATATTTCAAGTATTTACCAGAAAATTTGGCACTGGATACTACAGTGACTATAGAACCATCTTCAGTAACCTCAATGG tpg|BK006940.2|:62902-64414 24S84= 62=47S 
 tpg|BK006940.2| 105416 + tpg|BK006940.2| 105578 - INS TGAATCCAGCGGCACCGCCGCCGCCGAAGGCAGCGGGCCCAAATTGATCGTACTGCTGCCTCTTCGTTTCGTCTGACAGAATTTCATAAGCGTTCTGTAAATCGTGGAATTTCTTCTCAGCATCCGGTTCCTTGTTGATATCCGGGTGGTACTTCTTTGCCAGTTTGTAG tpg|BK006940.2|:105062-105932 11S104=19S 39S4=7X 
 tpg|BK006940.2| 151108 + tpg|BK006940.2| 151103 - INS CGCTTCTCAAACTATTACTTACAGACCCTTTTGTTAAGTGGGCTCTATGGATTGGCTATTGACTATACTTATACATTTAGTGAAATGGATGCGGTGCATTTGGCAATAGGGCTAGCAAGCTTGAAGCTATTTAAGATTGATAGCTCAACGCGCTTGACCAAAAAACCCAAAAGGGATATCAGGTTCGCAAACATACTAGCTAATTATACC tpg|BK006940.2|:150669-151542 7X111=46S 1=258S 
 tpg|BK006941.2| 221454 + tpg|BK006941.2| 221658 - INS TGTTGTATTCTTCCATAGAATATAACTCACGTTCATAGGCATGTTGTTCAACGTTCAATAATGAAGCCATTACGCCCTCGGAAGGTGCATTTCTAGTAACCTCGAGTAGCTCTTGAGTAATGGTTTTAAAACTTAAACTGTCAGTATTTTTTGGACCATTTGTACGTTCTATTACTCGCTTGAGTAAGGGTGTAGTAGAAACTCTAAAAAATTCATTCAACGAGGGTTCACCTGTTAATTTAGATAAAAA tpg|BK006941.2|:220940-222172 31S21=1X79= 102=30S 
 tpg|BK006940.2| 174303 + tpg|BK006940.2| 174482 - INS ATATTTGGATGATGCAGTCTTTGTAAAATGTCTAACTCGTCGTATAAAGCCTCTAGCTGAACCTTGTTTCCCTTTAGTGCTTTCTTGATCAGGATTTTAACGGCCACGTCCTCCCCTGTTTCAGTGTTTTTGGCTTGTCTCACCACACCAAATGTACCAGCACCTAATGTCTTCCCAAAAACATATTTTTTTTTATTCACGTACGAAGCAGGCTGCACATGTGCCATTTTACCTTCAGA tpg|BK006940.2|:173811-174974 7X5=114S 108S12=7X 
 tpg|BK006940.2| 37744 + tpg|BK006940.2| 37871 - INS AAACTGATGGTTCCGCTTCAATTTCACTTCCTAACCATATTCCATCTGTCAATCCTAGCAATAAACCAATCAAACGAATGCTAAGTAGCATTCTTGATATTAACGTTTCCTCATCAAAAAACAAGAAGTCTGAGGAGAACGAAATGATAAAACCCATGAACAAGGGCCAACACAAAAATAATACATCGTTAAACATAAACGGCTGGAAATTTGAATCTTTGCCATTAAAATCCGCCGAGAATTCAGGTAAACAGCAATATTATAGAGGATTGCCGTTATATGAAAAAAACACGCTGCTAGAA tpg|BK006940.2|:37126-38489 7X79=1X154= 151=7X 
 tpg|BK006940.2| 261336 + tpg|BK006940.2| 261569 - INS TTCTTGAGTCAAATTTTTTTGACGGAAACTTAGCGACCGAAAAATATATATGATAATAAGAAAACGAATGGCATACAATGATTAGTTTCAAATATTTCACGCGCAAAGAAAGAATTCTACTACCGGAGTGTGCCCTTCTTGTACTTTATTATCAGACTGTGTCTCTCTAATTGCGTGTTGTCCGCGGAATAATGCTCTAATTTAAAAAATCGACATATTCTGACTTGTATGGCGCTTTGCATTGGTG tpg|BK006940.2|:260828-262077 7X3=1I246= 124=7X 
 tpg|BK006940.2| 163659 + tpg|BK006940.2| 164408 - INS TTTTGGAGTATAGACGTACCCTGGGTCTACAAAAGATGCAATTATTATCCGGTGGTCAAAAATCTCGTGTAGCATTCGCTGCATTGTGTTTAAATAATCCACACATTTTGGTTCTGGATGAACCTTCTAACCATTTGGATACCACTGGTCTAGACGCTTTGGTAGAAGCCTTGAAAAATTTCAACGGTGGTGTCTTAATGGTTTCCCATGATATCTCTGTTATTGACTCTGTTTGTAAAGAGATTTGGGT tpg|BK006940.2|:163145-164922 7X9=10S 235=7X 
 tpg|BK006941.2| 981297 + tpg|BK006941.2| 980938 - INS AATTCCTTGTACCAATCAACCTTGATAACAGCTGCATCAAAGATATTTTTTGTTCCATGTCAAATTTGTTTTTCGTTTTGCCTGAAAGATGTTCCTTAAACAATTTTTCGGCAAATCCTTGTGGATCTCTCAAAAGGTGGATAGCACTGAAGTTTAAATACCCTTGAGGAGCACCCGGTCCGTTCTTCTTCTTCTTCTTCACAGTTTTTATGGCATTCTCCAGCTTCTTACCACGTCTACCCGTTTTTTTATTGACTTGCATCTTATGCCTTAATGC tpg|BK006941.2|:980370-981865 7X4=187S 260=7X 
 tpg|BK006941.2| 330223 + tpg|BK006941.2| 330513 - INS CCTGGACACTTCTATAAGTAAGTTCGAACGTTAACTAACTGTAATGACGTTACCCTTTCCTGAAATTGGCAGAAACAAAAATGAACATTTCTGGCAACTTTTCGCCATACAGTCAGTACTCGTTACGGACGCCCGGGAAACAAGTAGGAAACATATGAGAGGCCAAACAAGGGTAAGACCTTCTTTTCTGGTAATAGATATTACTTCAT tpg|BK006941.2|:329791-330945 7X191= 105=7X 
 tpg|BK006940.2| 109755 + tpg|BK006940.2| 110513 - INS ACATTATGTGTAATGGAACTCGTATCACACATTGTCATTGAAATAAATCATTCACCTACCGCAACAACGGATGAAACGAGAAAGCAGAATAATCCGGAGCTGAAAGTGAAAGAACCAGTTTGTAACCTCAAGAAGTGGGAAAATAACACTAACTTTATATTGGAAGATCATACGAAGAATAAAACAAAACTTTCTAGCACAGATAGGATACGTAAG tpg|BK006940.2|:109309-110959 7X194= 203=7X 
 tpg|BK006938.2| 830658 + tpg|BK006938.2| 830760 - INS TGTCTTGTCTAGGATAACAATTGAATACAAGATCTCGCGTAACCTTCTTTAATAAAATTGAAATTGAGCAGCAATTTATGAGTATTAATTATTCTTGCCTTCATTTCCGAAATTTGACTTATTGTAAACTCATTTGTGAACTTAGCAGGCTTCGTTGCAGATACAATGTCTTGTCTTGCAGAATCTATTTTAGATGTTATATCAGTAATCATGGATTCTATTTTTAGGTGGGATTCATTAGCGTCGGATGAAGCTAACGAAGATGAAGGTGATAGGGATGCAGGGGATAACATGGGTTCATTTGTGGTTTTCAAAAGGGATTTTTTCTTCTTGATGGTGGGTTTATCTATCTTATAGTTCTTTTGTTCTTTATCAGGTTTATGTACGTTATTTTGGTTTGTACTTTTATCTAATGATGCCTTGCCAGTATAACCCTTTTTATGCCTATCGAGATCAATACCAACT tpg|BK006938.2|:829714-831704 7X304= 3S448=7X 
 tpg|BK006941.2| 985252 + tpg|BK006941.2| 985951 - INS CATACATCCACAACCACCTCAAGAAAAATGGTGAAATTACAAAGGTTTAGCGAAAAGAAAAGCCTCATACACGAATTCGGCAAGTTTATCCTTGAAAAGCAAGAATCGGCGTTAACGGGCGACGCTGATGCAGTGTTCAATATCGCCATCAGTGGAGGATCGATGAACCAAGCGCTGTACGAAAGTTTGGTAAATGACAAAAACATTTTTCCACATATTAAGTGGCCACAATGGAGAATCTTCTTCTGTGACGAAAGATTGGTTCCATTTGAGGATCCGCAAAGTAACTATGGTCAGTTCAAAAAAACAGTTTTGGACCCGCTAGTGCATCAGGGCAACCAATTGAACTTAGGCCCCACTGTATACAC tpg|BK006941.2|:984502-986701 7X169= 184=7X 
 tpg|BK006940.2| 71701 + tpg|BK006940.2| 72125 - INS TCTACGGAAGGTTGAGGTTGAAGAGAATCTTTATCTCTAGACAGCATTTCGTTGGTGCGGTCATCATTATCTACATGTGAGTATTCTATCTTTTGTCTTGGTGTTATGGATCTTGATCTTATCCCCAGCCTTGACGAAGAGGAAGAAGGTCTTTCCGAGTTACTAGTCCGAGAGTCGGTGGCTTCACCAATACCATACTGTTTCATACTACTACCCCTACTA tpg|BK006940.2|:71243-72583 7X159=35S 23S5=7X 
 tpg|BK006938.2| 205724 + tpg|BK006938.2| 205869 - INS TTCTTCCTTCTCTTGCTTTGGAGACGTGGCTTCACCATAATCAGCACCACCGTACGCTGTAAATCCTCCAGCCATAGCGTCATTTGAACCCGAATCAACCAGAGGTGAAAACATTAGCTCATCTTTAACGTCAAGATCTGCATTGACCAAACCACTTTCGTTACTGTATGGTGTGACGCCACCATCTTGTCCGTCTTCAATCTCAGTTATTTTTTGTTCTGGCATGTATTTTACCAGTGACTCCTCATCGATCATCACATCAAATGCACCGGTAC tpg|BK006938.2|:205160-206433 7X179= 1S257=7X 
 tpg|BK006941.2| 594103 + tpg|BK006941.2| 594046 - INS TGGTTACATACCACCATATTTTATCTGATGTTCGGCGATTGCCTTTTTAGAGTCTCCAAATCAAAGAAGGTTCAGCATCTAAAAAATTTCGATGAGTTTGAAAAAGATCCATTTGCATTCATTTACAGGAAATACGTAGTACCAAGGCTCTCCTGTGGTTACAATGA tpg|BK006941.2|:593698-594451 183S68= 147=7X 
 tpg|BK006941.2| 2363 + tpg|BK006941.2| 2580 - INS TCATTACAAATACTCCGGGTATAGACACTGAAGACTGGGAACGTGTTGCAGTAAATTTCAATTCTTATTTATATGAAAATAAACTTTGGAATACTGAGTACTTTTTTTTTGATGGTTCCAGCTGCCAAGAAGCGTTCAGAAAGATGCTTCTTGAGCCATTTTCCTTGAAAAAAAATGACTTTGCTAATGCCAAGGTACCTGACGGATCTGTTTGTTAC tpg|BK006941.2|:1913-3030 7X6=103S 101S8=7X 
 tpg|BK006941.2| 7208 + tpg|BK006941.2| 7338 - INS CCCATACTCATTCCCAGAGGAAACACTTTGCAGTAAGAAATCTTTCATTCCCAGAGAGAACGCGGAAATATTCAGCCTAAGTCTCTCCAAATTGATTTCTTTCATTTTGGTAGCGAAAGACTTAGTATCAACCTCAAAAAGCTGAAATTTTTGTAGATATATGTGCAGATGACATGAAGTATCCAGCTCTTTTGTGAATATGGAAGCAAGTTTCTTTCAAATTATTATCGACTTTTCCTCTGCCCCTTTTACCTTATAACTTTAGGAAACACTACCCTATTC tpg|BK006941.2|:6630-7916 114S60= 2S5=1X257=7X 
 tpg|BK006940.2| 190999 + tpg|BK006940.2| 191508 - INS GTGGAGGAACTACGCAAACCGGGGATCCTTCTGTTAACATTTCTCCCTCAGTTTCTACAACTTCTCATAATAAGGGGAGGGACTCAGAAATTTCATCCTTAGTAACCACCAAAGAGGGCTTGTTGAACACCCCTCCCATTGAAGGCGCCCGAGATAGGACCCCACAAGAATCACAAACGCATTCCCAAGCAAATTTAGATACTCTTCAAGAATTAGAGAAAATTATGACAAAAAAAACAGCCACACACTTGAGATAT tpg|BK006940.2|:190471-192036 7X4=124S 114S15=7X 
 tpg|BK006940.2| 26823 + tpg|BK006940.2| 26623 - INS TCTATATCTCTTGAGCGCCAATATGCGAAAGCTTTCACAAGGTTGATGTTCATGGTATTCGGCGTCGATAGCGAATTGCTTACTAAGAAACATTAGGGTGCAGTACAGCCTTGTTTTTCCAGTTCGACTAACCTTTTTCTTGGCAGTATGGAGAC tpg|BK006940.2|:26299-27147 7X40=37S 1=158S 
 tpg|BK006940.2| 82243 + tpg|BK006940.2| 82162 - INS GTTCTCTTATTTGACTTCAAAGCAATACGATACCTTTTCTTTTCACCTGCTCTGGCTATAATTATAATTGGTTACTTAAAAATGCACCGTTAAGAACCATATCCAAGAATCAAAAATGTCTGATGCGGCTCCTTCATTGAGCAATCTATTTTATGATCCAACGTATAATCC tpg|BK006940.2|:81806-82599 11S131=16S 15S5=7X 
 tpg|BK006941.2| 618819 + tpg|BK006941.2| 619217 - INS CTTCATCTCTCACTTCATATGGCAAGTCATGCCTTAAATTGTGAGGATGAGGTTCTACAGCTGTAGTTTCTGCCGTAACGTCTGTCTTCGAGGACTTATCTACGCTATGATGTAGCTCCTCTTCAGCTATGATACTGGAGTTAGTATCGTCTGAGTATAAG tpg|BK006941.2|:618483-619553 7X6=74S 76S5=7X 
 tpg|BK006941.2| 494438 + tpg|BK006941.2| 494578 - INS GCGATCTATACTGCTCTCTGAGCCTACCGTATCCTTGCTTAGCATCTCGCCAAAAAGCTCATTCTTCAGCAAAGTATTATAAGTTTCATGTGCCTGTCTTTCCTTTTGGTATTCTACTTGATCTTCCGTACTCGATGGATTAAGGGCTGGAACG tpg|BK006941.2|:494116-494900 7X3=74S 73S4=7X 
 tpg|BK006940.2| 249921 + tpg|BK006940.2| 250185 - INS GAGTATTTAAGGGAGCTCTTAATGGAGGTTCCCATTTCTTGGTCCATGTTGACAACTTCAGCGTCAGAGCATGTAGAAGACTCTGTATTTATGTCTACTGGCTCCTGAGGGAAAACTGGAATGGTGAAGATCACATCAGCGAGTTCTGTTTCCAGGACGCTCTCATACTCAATAATGACATCAAAGCCCTGTTGTGATTCGGAGGGGGAAACCCATGTAGTTAGAGTTAATGGAATTAATG tpg|BK006940.2|:249425-250681 7X17=1X32= 1S225=7X 
 tpg|BK006940.2| 207495 + tpg|BK006940.2| 207983 - INS TACCACCTTTATGGGGGCAATGGTAAAACATCTAGTCGTGGACGTTGGATGGTTTATGATTCTAGAAGATTGGTACAGAATGTGTACCCCGATTTTAAGATTGGCATATCGAGAATTTGGGTGTGCAGGACAGCAAGGAAGTTGGGTATCGCAACCAAATTGATTGACGTTGCAAGAGAAAATATTGTTTACGGTGAAGTTATTCCTGGGTACCAGGT tpg|BK006940.2|:207045-208433 7X223= 98=1X10=7X 
 tpg|BK006940.2| 147549 + tpg|BK006940.2| 147296 - INS ACTATAACCTCCAGCACATCGAGGATAACAAAAAGCGCAAAATTTCGCAAGAAGAGGTTACGAGAAGCAAGGCGAAAAAGGCTCCGAAGAAGTTTGACTTTTCTAAACATAATACCAGGTTCATCGCCTTGAGATTTGCCTATTTGGGATGGAATTACAATGGCTTAGCTGTTCAGAAGGAATACACACC tpg|BK006940.2|:146902-147943 7X5=220S 167=7X 
 tpg|BK006940.2| 96117 + tpg|BK006940.2| 96386 - INS TATATATATATTCCTCCGTGAGGAAGAAGAAACCTGCTTTGAAGAAGATCAAGTCTTCCACTTCTGTGCAATCTTCGGCTACTCCGCCTTCGAACACCTCATCCAATCCGGATATAAAATGCTCCAACTGCACAACCTCCACCACTCCGCTGTGGAGGAA tpg|BK006940.2|:95783-96720 7X11=69S 77S3=7X 
 tpg|BK006941.2| 965317 + tpg|BK006941.2| 965322 - INS CTAAAATCCCCCTAGAAAAGCGGGCTCTTTACCCGGCGAATAATAATAACCGCGGCTACTAATTTTGCACCATTGAATATTAACCTCAAAAGGCTTAGTTGGCAATTATATTCTCCTTCTATTAATACTTAATGTTTACAATGTCCTTATAGGTGTTTAAATATATTTTTATATACTTTGTAC tpg|BK006941.2|:964937-965702 7X3=88S 89S3=7X 
 tpg|BK006938.2| 1033690 + tpg|BK006938.2| 1033285 - INS GGATAAGCGGATGAAATGGGAGTACAAGAAGAACTATTAACGTCATCAGGGAATATTCAAACTGCTTTGGTAAGTGAAATGAATAACACAAGGCAAGAGCTTCTTGATGATGCGTCTCAAACAGCCAAAAATTACGCGAGTTTGGAAAACTTGGTGAAGGCATATAAGGCAGAAATAGTTCAGTCGAATGAGTATGAAGAAAGGATAAAACATTTGGAGAGTGAAAGGTCAACTTTGTCTTCACAAAAAAATCAGATTATTAGCTCTCTTGGTACTAAAG tpg|BK006938.2|:1032711-1034264 7X163= 263=7X 
 tpg|BK006940.2| 134048 + tpg|BK006940.2| 134641 - INS CTATCTACTGGTCTTTTGATCAACAACGCCATTTGAATCTTCGTTTTCAGTCCTTGCTTTTGCAATTTTCAAAAGCGAATGGATATTGTACGCTTCTGCAATAATATCCGGGTTGAATATTTTTTCTACCACCCTTATTCCACTATTC tpg|BK006940.2|:133738-134951 7X10=146S 107=1X22=7X 
 tpg|BK006941.2| 12411 + tpg|BK006941.2| 12312 - INS GTGCAATTTTGGAACATATCATTTAGTCTCTGTCTATGCTCATAATCGTATTCCCATGAAGTTTTTTTACAAATATTAAGGCCCCCGTTTAGCCATAGCAAGGACCCGTCCCTGTCTGTATGAGATAGTTGCACAGAACAAATCTGGTAAAACTCACCGGTACTCTCTTTTGAAACTACATTGCC tpg|BK006941.2|:11928-12795 12S96=37S 42S5=7X 
 tpg|BK006941.2| 863084 + tpg|BK006941.2| 863321 - INS ATAGACCCAAAACCCGACGTCAATTTGAGAGCACAATACAACTGATCTCAAAGAGAAATCCGATATTTTCAGAAAATCTGAACAGTCTTCTAACGCTTCGTATGCATCCTTTAAAGACACTTTTTCGATAAGGAATGAAAGCATTGTTTGTAAAGGATTCATAAATGCAACTCTTTCGTGGCTTACGCTAAACTTAATGACTTCATGAGAATCATATATTAACTTGTATGTTAGTGATCTATTGCCTAGAAATGAACTGATAATTC tpg|BK006941.2|:862538-863867 7X245= 133=7X 
 tpg|BK006941.2| 125109 + tpg|BK006941.2| 125616 - INS TGTTTGGAAATCGCATCATCAGACGATTTTGTTGGGTACCAAGACTGATGATTATTATTCACCCAGTGTACAAAGATTCGACCATCTTTCCACTTTTGGATTACCGCTGGTAAATATTTTTAACAAGACGATCCAATTACCCCATCACAAGATCTCAGCTTCGTCTTTACCAATACCCATAGAAAATTTTGCGAAGCATAAGGATACTC tpg|BK006941.2|:124677-126048 7X92=64S 2S1=303S 
 tpg|BK006940.2| 260742 + tpg|BK006940.2| 260875 - INS GGAATGTTCTTCTGAATCTGAATAAGGTCACTTACATAGAAACCTACTTACCTCAAAAGCGTAATTCCGAAAGGCAAAAGAAAAACTTTTGTAGAATCTTCAGCTGCTAGAAGTTCAAATAGAAGACAAATTACGGACTTGTTGCAGTATATGCCAAGCTACAGAAGAAATTATATTTCTTAATACGTACAGAAGG tpg|BK006940.2|:260336-261281 7X7=7S 98=7X 
 tpg|BK006940.2| 193842 + tpg|BK006940.2| 193748 - INS GATCTTCTTGTTCGTGGGCACACTTACTTAGATATTTCCTTGCGCAGTTATTATACTGAATTTAGAGAAGCGACGCAATATTTCTACGTGATATCTATAAAAAAGAATACTTCACTTATGCAAGCATCGCCTGGCTGTAATCTTTGCTTCAGACCATCTGACACATGTACAC tpg|BK006940.2|:193390-194200 7X6=265S 86=7X 
 tpg|BK006941.2| 471156 + tpg|BK006941.2| 471303 - INS TTGACATCACAGTTGTATGTCAAAGTTGCCTGTGATTCGCTATCGTCTTCATAAAAACCGTTTCTATTCACATCGTCGTCATTCTTCCCATCACTTCCGCTATTATCACCACTACTACGACCACCTAGCTTGAAATTCTCAAAAAATTTCGTTGGTTGTTCCACTGCGCATGGCCCGTCTGTACATCGCTGAGGATTAGAAAAAGAAGTCGAACTGGAATCTGTTTCCTCTTTGACTTGTACGGTTGTACCTTCCAAACTCGTCTTGTGAAGGTTTTTTATTCGAGCGCCACCTTGTCTAGTGC tpg|BK006941.2|:470534-471925 23S136= 148S4=7X 
 tpg|BK006940.2| 252421 + tpg|BK006940.2| 252019 - INS GCTATTCAAGTGATGAGGCGGAAACGTGCAAGATCCTAAATGAAGGATAAAAAGAGTTCTTAAAAAGGGAAGTAAGGAATAACAGAGTAGAAAAACCGAAAAGACAACTTAACAAATCGGCAACACTTTTATGGGGCCCCGCTCGCCTGTGTGCAAGTAGTATTCGACCTGGAACACGCATTTACCACGAGAAGACAGCAATAGTCCGTACAACATTAATTAGTTTCGACAATTGCTCGCCTTTATAAGCCATGCTAGTGCCCAATCAAACACTTTACTTGCCCTGAAGTTCCTTTTTTCGCTAGCCTGTAACTTAAATAAGCCATCTAACCTTTTTTTTCTAAAAATTTTCTTTATTACCCTGTCGGCTTATTTTCTATTCTACACATTATTTGCCACCCATTGAAATTGTAGCT tpg|BK006940.2|:251173-253267 7X5=106S 208=7X 
 tpg|BK006941.2| 737172 + tpg|BK006941.2| 737681 - INS TGATTACCTCTCTAGGTTGGCTGTTCAAATTCTAACTTTGGACCTTCATAATTGGCTAAATCTGCATTAGCATCAAATGAACTCAAGTTCAAAGTCTGACACAAACTGATCTTGGCTTCATTTTCTGCGCCTCCGATAGCTTTCCTAAATCTTTCTTCTCTAATGAACCTATCACATGTAAGTAACGCCTTAGTAGCAGCCGGATCATTGGGCTTCGCCTTTAGAAGCACATTCAAATCTTTCCTAGCCTTTTTAAATTC tpg|BK006941.2|:736638-738215 9S246= 3S241=7X 
 tpg|BK006940.2| 244238 + tpg|BK006940.2| 243904 - INS TCTTCAGATTTGTTCTTAAGACTTTGGGCGCACATTTTCAAACCGTCACCTTTGAAATTATCCAACATGATAACGTCTGCACCAGCTTCAATGGCCTCTGTGGCTTCATCTTCACTCAAACACTCCACTTCGATCTTCACAGCAAACCCGCACACGGCCCTGGCG tpg|BK006940.2|:243560-244582 14S137= 14S7=7X 
 tpg|BK006940.2| 158520 + tpg|BK006940.2| 158441 - INS AAATGTGTACATAAAAGTGGAGAAACAGTTATCAACCCTAATGGAAGCTGAAATGCAAGATTGATAATGTAATAGCATAATGAAACATATAAAACGGAATGGGGAATAATCGTAATATTATTATGTAGAACTACCGATTCCATTTTGAGGATTCCTACATCCTCGAGGAGACTTCTAGCATATTCTGTGTACATAATATTATGG tpg|BK006940.2|:158019-158942 7X4=173S 6=1X185=7X 
 tpg|BK006940.2| 21362 + tpg|BK006940.2| 21718 - INS CCCTCCCGAGAAACTCCGCAAACGGTTCTCGCATATGATAGCGAATTTTTGCCCAAAAGTTAGGAAATGTCATTATATCCGCGTCTTCATCTTCTGAGGCACCAATTTCATTACCATCTAATGCACTCGTACTTTTATTTTCCTCTTCAATAAGTTCTTCAGGAAGCTTCGTATAAACCGGAGTAGAACCATCGAGGGTTTGCATGTTCTTTAATTTTCTGGATTCTGCATCGGCTATGGAGGA tpg|BK006940.2|:20860-22220 7X5=12S 122=7X 
 tpg|BK006938.2| 934299 + tpg|BK006938.2| 934765 - INS TGTCATTTATTAAAAGGTATAAATATGTAAATGTATACTTAATGACCGTTAAGAAAAACTACTAGCCTCATCACTCCCGCAGATCTCTATAATTGTTGTTTGAATACTTGATACGGTGGAGTGGCAAGGACAGTCTGCGCAGTCCTAATATCGATATTGATGTCTTCGATCAGAGCTTCCTTAGTAGTGTAGTTCAATTCGGGTCTGATATGACCTAAAATATTGAACTTGACCCTGGCCCCATAAAAATCATTTTTAAAATCATGTATAATATGTAATTC tpg|BK006938.2|:933723-935341 7X192=18S 1=159S 
 tpg|BK006940.2| 103119 + tpg|BK006940.2| 103518 - INS CGCATATAGAGTATTGCTGAATATAAATGGATCTAGGAAAGTGGCAGGAATTTTGCGAGGCTACGATATTTTCTTAAACGTCGTTCTTGATGATGCAATGGAGATAAATGGTGAAGACCCTGCCAATAACCACCAGCTAGGCTTGCAGACCGTCATTAGGGGCAACTCCATAATATCCCTAGAGGCTCTAGATGCCATATAAAATTATATATATATATATATATGTCGACCTCTATGTACTAT tpg|BK006940.2|:102619-104018 7X145= 228=7X 
 tpg|BK006940.2| 81196 + tpg|BK006940.2| 80929 - INS CTGGTGTAATGCACC tpg|BK006940.2|:80885-81240 7X4=3S 3S5=7X 
 tpg|BK006941.2| 630833 + tpg|BK006941.2| 630569 - INS GGATCTCTGTTCAAAGACGGTTCAAAGACCTATGCTTTTAAATCTACATGATAACAAAGTTTTAGCGAACATGTATAAAGAGACGTTCAAAGTAGTTTCCATGTTTCCGATAAAAAATTCAACTTTTGCATGTTTTCCAGAACTCTGCTTTTTTCTCAATAAGCAAGGGAAGAGGGAGGAGACAAAGGGATGTTTTCATTGGGAGGGGGAACCAGAACAGTTCGCGTGTTCCTACCCTTATATTGTGGCAATTAATAGTAACTTTATTGAAATTAGACATATAGAAAATGGAGAACTTGTCCGCTGTGTACTTGGAAACAAGATACGTATGTTAAAATCATATGCCAAGAAGATCTTATATTGTTATGAGGATCCTCAAGGATTTGAAATTATCGAACTGTTAAATTTTTGAGTTGACCGCCCATATTAATACCTTAAAACTTATTTCTTGAACCTATAC tpg|BK006941.2|:629635-631767 13S7=1X145= 5S427=7X 
 tpg|BK006940.2| 258056 + tpg|BK006940.2| 258197 - INS TAGGTGAATGACGATAGAC tpg|BK006940.2|:258004-258249 7X4=5S 10=7X 
 tpg|BK006941.2| 421935 + tpg|BK006941.2| 422131 - INS ATATAAATGTAAAAGAAAATAGGAATTGCTGTCGATAGATTTATTTACTTTTGTATTGTCATCTGTGTTCTGTGCCAGTACACCGGACTCGTATGAGCTGTATGGTGTCGTTTCAATAGAATCTACTGTAATAATCACACAGATTAGAAATTATTTTC tpg|BK006941.2|:421605-422461 7X7=72S 73S6=7X 
 tpg|BK006941.2| 748879 + tpg|BK006941.2| 748938 - INS GGACAAGAGTTGAAATAGCTGCGTGCTTTGGCTAGGGTTGAAGCATTCTGGTGAGCTGTCTTCACCACCGCTTGTTATGAACTCAATGAAATTTTGAACGTCTAATTTACTTAGTTTCTTCATTTCTTGTTTAATAGAGTCTCTGGTGAAATCCTGCAAAAT tpg|BK006941.2|:748541-749276 7X4=77S 76S5=7X 
 tpg|BK006941.2| 981719 + tpg|BK006941.2| 982326 - INS TGACAATCTTAACATCCTGATGTAATGCTGCTTGGGTCATAATTTCTACTGTTCTTGAATCATCCCAAATACCACGTCTCCAAAGTTCTCTGGTTAATTTTGTGGCCCAGATTCCCTGGGAATCTGGTTGATCTAACAAATTAAAGCAAACGGCCTGCGTAGATTTGTTCAATTTTTGATTTTTACCATTAGTATTACAA tpg|BK006941.2|:981305-982740 7X3=281S 100=7X 
 tpg|BK006941.2| 422943 + tpg|BK006941.2| 422986 - INS AACAGAAAGTTCCAATGGTTATCTATAGGTTCCGTTTCAGCTTTACGTACCTCCCAGTCAAGGTACGATTCAAAGCCTTTTAATTTTTTATCCCAAATAGAGCACGATGTCGCAATCTTCTGAGTGTTAAACTGTCGCCAAATCTGTATTTGGGTATAGCCATTTCTTCCAAAATTGCTAGGAATGGCCTTATAAGCTATATTGTGCTTGTGCTT tpg|BK006941.2|:422499-423430 7X7=100S 102S6=7X 
 tpg|BK006938.2| 845704 + tpg|BK006938.2| 845516 - INS GCGTAGAGGAGGAAGAGTAGGATCTTCGAAAATACAGGCGTCTTAATAGAGGAATTGTTATTTAAAATACAACCCACATCTCTTGGTCCTCCTTTTTTATCTTTTCTAATATATGTTGCTGTTTCTACTGGAGTAATTATTTTTATCATTACTACGGGAGAATGAGCGTCTATTGTTGTTGCTGCGTCTAAACGGTTCGTCATCGTAATCTCTATTTTGGCTCCTATTATTATAGTTTTTGTTGCCTCTGAAAGAAATTTCTGAATCATCATCATAATCGTAGGACTTGTTATTTCCATCTCTACTACTATAGTC tpg|BK006938.2|:844872-846348 7X288= 9S287=7X 
 tpg|BK006938.2| 856115 + tpg|BK006938.2| 856282 - INS ATGGGTCAAGAATACGAAGGCAGAGACGCGGACGACGTGGTTATGATGGCATCTTCTACTAATGAGGAATTGGAAGAATTGAAGAAACTAAAGGAAAAGAAGAAGCAACTGGAGAATAAGTTGGAAATACTCAAACAGAAATAGTTAGAAGTTTATTTTTTAAAGCATCCATTTATCTCTTTATCCAGTTTGTATTATAAATTATTGTTAATGTTATCGCTAGTAGATTACTTATATGTACTTAACTGTTTGCTAGCTACCAAATTTGCTTGATGGTTCGCCATCGAAGCTTTGAGACTGTTCAATTTGGCGCTTATAC tpg|BK006938.2|:855463-856934 7X264=15S 1S1=236S 
 tpg|BK006941.2| 621466 + tpg|BK006941.2| 621555 - INS TACATCATTTTTCCCTACTTTCTTTTTCTGTAATGGTTCATCGAAGCATTTTTAAGGGTGCCCTGAAGACTATTGTTAAAAAAAGGTACCGCATACATTCGAACCATTACCAGAAAAAAGAGGGGTGAAAAGACATTCTAAATTTTGTTATCGAATGTGAACAGAACACTTAAGAAAACGCCAAGGTTAAGAAGGCCTTGAGAGTATTGATTAAGGCGCATGGAGCACAGGTAAACGCGAAAGACGTTTTGTACTTCCTTTTACTGAGCACCTCTTACATGTAGTAG tpg|BK006941.2|:620878-622143 7X214=37S 17S1=239S 
 tpg|BK006941.2| 729199 + tpg|BK006941.2| 729121 - INS ATTTCAGTGGATCCCGAAAAGTATTTGTGGCCTGATTTGCACCAAACCCTCCGGTAGTAGCCGTCCCAGAATTTGGCTGGCTGCCCCCAAAACCAAATCCTGAAGCCGAAGGTTGAGTATTTGTATTGTTATTGTTTTGTCCAAATGAAAAACCGGTCGAACCAGCTGGTTTATTTCCGAACCCGTTATTACTACCGCTGAAACCAAACATGTGATCAATTGGTCAACAAGGTATGTC tpg|BK006941.2|:728631-729689 23S103= 110=16S 
 tpg|BK006941.2| 867646 + tpg|BK006941.2| 867633 - INS AATGAGAAGAAATTTCCTGAGGATGAGAATGGGTCAAAACGGCAGCAATTCTAGTTCCCCAGGCGTACCAAATGGAGACAACAGCAGGGGATCTCTTGTCAAAAAGGATGATCCTGAGTATGCTGAAGAGAGAGAGAAAATGCTTTTGCAAATCGGTGTCGAGGCCGATGCTGGCAGGAGCAATGT tpg|BK006941.2|:867247-868032 7X93= 155S3=7X 
 tpg|BK006941.2| 164173 + tpg|BK006941.2| 163926 - INS GTTATTGACATAGCAACGCCAAAATCGGATATTTTCACCGTTCCGTTTGATGAAATTAACAGGTTCGATGGTTTGATATCTCGATGCGTTATCCCTTGGGAATGTAAATACTCCAGACCCGATACTACATCCAACACTACCTTCCTCGACTGTTGGAAAGTGAGTATTGATGGTCCCACTGCTTTTATCTCCATTTTGTTTTCTGGACACCATTTAACGGGTCCCCTTGAGC tpg|BK006941.2|:163448-164651 11S200=13S 10S5=7X 
 tpg|BK006941.2| 615312 + tpg|BK006941.2| 614965 - INS GTAGAGGTCCAATCAGCATTGAAGATCGTGTGACGACAATGTTCAGAATTAACTTGAGCGAACATAAATAACTCAACATCAGTAGGATCTCTTTTCATAGTTTCGACGAATGCATGAATCAAATATTCCATTTCTCCACTATCTAGAGCTAAACCCAATTCCGTATTAGCTTTGGATAAAATATCCTTTGGAGACTGTTTAGTGT tpg|BK006941.2|:614541-615736 7X4=208S 103=7X 
 tpg|BK006938.2| 1490899 + tpg|BK006938.2| 1491225 - INS AAGTGATGGAAGGAAAGACTAAGAGAAAAAAGAGCCCAAAAGAAAAAAACTAGTGGCAAGGATGCTGAAAAGCAACAAACGAGTACAGACGCCCCACTATCCGAGGCAAAATCTATCCATAATGAAAATATTAAAGTTCTGCAGGGAATGAGTGATGAACAAATCGTGCAAGAACGTGAGGATCTGTATAACTCTTTAGATCCCAAACTGATTGCCAAGCTATTGAAAAACATAAATAAAAGAGCGAAGGACGAAAACAACACTCCATTATTTGCAGAAATAGAAGGCGCTTCTGGTACCTGGGTAGGTGGCAACAAGCAAGGCATATAC tpg|BK006938.2|:1490225-1491899 7X149= 165=7X 
 tpg|BK006941.2| 132360 + tpg|BK006941.2| 132724 - INS TTTTTGAGTTATGCTGCCTCTGCAAAGGGCTGTCCCCATATATTGGTAAAGAAGGTAATGAAGCAGCCTTGACTCTAATGCTTAACGCTTTTTTTGTTCATTATTTTAGTCTGGGCAAACCTATTGAAGACTTGGATAAAATTATATCAGCTGGTTTTGCAGATAAAAAACCTGCTTTGAAAAAATGCTGGTTTGCCGCATTTTTGAACAATTCCAATGCTGCCTCTGAAGAGGTGATTTTAAACTTTATAGACGGTTGTTTGGAATTTGTGAAAGACTCCATCATACATTATCAGACTCACGGGCATGCATGTATTCTAGCATCAATTGAATTTACAAACAAAATTTTGGCATTGGACAATACTGAGCTAAATGATCGTGTTATGCAGCTCATAGAAACCCTTCCTGAAAATTCTTCGATAGGTGATGCTATCTTAAC tpg|BK006941.2|:131468-133616 7X6=102S 5S421=7X 
 tpg|BK006941.2| 276964 + tpg|BK006941.2| 276327 - INS CCATTGACTTGAAGAATGTTTCATCTAGATTAACCGATGTCGTTGGTTCTGAAGTCGTTGCCACGATTGGAATACCCTCAAAATTCCCACTTTTACTATGCTTCAATTGACCCTTCGGTATCTCAGCATCTAGGTAGCTTTCATTGAGATTCATAGTTCCGATGTACTGATTCTACGTTTGTGT tpg|BK006941.2|:275945-277346 7X10=148S 92=7X 
 tpg|BK006938.2| 1290225 + tpg|BK006938.2| 1290987 - INS GGTAGAACTTAATAATAATAATAATAATAACAATAATAATAATAATGATAATAATAATAGTATCGAAAATAATGATAGTAATAGTAATAATAAACATGATCATGGTAGTCGCAGTAATACTCCCAGTCATAATCATACTAAAAATTTAATGAACGATAATGATGACGATGATGATGATCGACTTATGGCGGAAATAACTAGCAATCACCTTAAAAGTACTAATACAGATATTCTAACTGAAAAAGGTTCAAGTGCACCCTCGAGAACCCTGGATCCAAAAAGTTATAACATAGTTGCTTCAGAAACTACTACTCCGGTGACAAACAGGGTTATTCCTGAGTACCTCGGAAACAGTTCCAGTT tpg|BK006938.2|:1289487-1291725 7X216= 340=7X 
 tpg|BK006941.2| 174698 + tpg|BK006941.2| 174695 - INS AAGAAAAATCAAACTGCCTCGAGTCTGACGATAGAAGACCCTGCAATAACATTTACACATGACAAAGAAAGAACTGTAAAAACATCTTTACTGGGCCGCAAGCTTTATGATAAGCCAGCACCTGAGAACAGGTTTGCCATTATGCCTGGGTCAAGATGGGACGGTGTCCAC tpg|BK006941.2|:174339-175054 7X7=78S 82S4=7X 
 tpg|BK006941.2| 382321 + tpg|BK006941.2| 382866 - INS TATGAGTTTATTCGTATTTGTCTATGAAAGGTTTCACAGCGTCTCTGACAGGTGGAAGTATAAGCAATTGGTCGAAATTCGATATTTTTTGAATGAGTTTATTCGTACTGTCCATATTCATCTCGACGTCTTTTTTCAATCCACCATACTCTCCAAAGTTGAATGCTTGGTCAGGGTCATTCTTTTTGTTACCTTTTTTGCCTTTGGCCTTCTGTTTTCGGTTTTTATTACTACTGCCTGTAGGCACTGAAGCTAATGGAGAGTTTCCTTTATGCTTTGTTCTTGGGCCTCCCGCATAAGAACGCACTCCTATCTTGAGAAGCACGGGGAAAGACCACTGTGGTGAAATTACTGGCTTGAAAAAAAGCGACATTTGTCTTATTATACTTTAATCTGATCTGAAGAAGTATTTCTACTC tpg|BK006941.2|:381471-383716 7X174= 66S326=7X 
 tpg|BK006938.2| 1131689 + tpg|BK006938.2| 1131586 - INS GGCGTTCAGATAAAAGAGCTTTGTCAATGGTAATGGATAAAATTGTGTACCACCGGGGAATACTGGAAATGATCGATGACAAGTGGCTATGTGAGGCAAAATTCACGTCAGTCAAAATTGAAGCAGACTTATCAGATGTAAAAAGCACTGCAGATGACTTCCAGCTGGCACCGTTATCGTCTCTAATGAATACGAAAGAAATTAATGAAGTAATTCTGAAAACTTACCTTCATAAAAAGCAAGAGAAATCACTAAAATCAACATTACTGTTTGGCGTTGATAAAGCCCATGTACAAAGTTTGCATAAATTATTTAAAGACAACGGTATTAATA tpg|BK006938.2|:1130906-1132369 7X178= 167=7X 
 tpg|BK006941.2| 59209 + tpg|BK006941.2| 59567 - INS CAATTCTATACAAATGTATGTTAATAACAAAAAAATTTCACTAAAAATTTCAGAAGCAACAATTTTAATCACTAAGGTTGTTAGAATCTTGGAATTATCCAGCAAATGTCAAGAATTGATCACCGAAAGAAAGTTTTTCAAAGTTTTACAAAACTTGGATAGTCT tpg|BK006941.2|:58865-59911 7X11=145S 145=7X 
 tpg|BK006941.2| 316623 + tpg|BK006941.2| 316086 - INS ATAGGAGAGTATATATTGAAAGATTACGTCAATGGGAAATTACTGTATGTCAACCCTCCGCCCCATCTAGAGGATGATACACCTCACACTAGAGAAGAGTGTGAAGAATTTAACAAAGATTTATATGTGTTCGACAGATTACCGGACACCAGAAAGGAGCAAGTGCAAAATGCTGCTAAGGCTAAAGGCATTGATATCGTGGATTTAGCTCGTGATTTGAATCAGCTAACGTTTTCAGCTCACACTGGTGGTGACACACAAAAAGAAGCCAAATCTGTTACGCACGGTGGTAAAC tpg|BK006941.2|:315482-317227 7X5=394S 66=1X210=7X 
 tpg|BK006941.2| 67153 + tpg|BK006941.2| 67451 - INS AAACGCTTTGCCATTATACCAATCCAAGAGTCTGGAACACCTACTTTTCAAGAAATTGTGAATTATACAAAAATAAAGTTAGTCCCGGTTTCGATATAGTGGCGCGTAAATATGACACGGCTGTCAAACCTGTCATCGATGACGCTACAGTAAAAGTGAACAAGGTCGCTATACAGCCTGCATTCAAGGTCATCCATTCACAATGTAAGAAATGGAACTGTGGAAAGT tpg|BK006941.2|:66683-67921 7X114= 232S4=7X 
 tpg|BK006938.2| 1051900 + tpg|BK006938.2| 1052071 - INS ATCATATTATAACCATGGGGTATTTCTGAGGTAACCATGTATGGCTATTTTTAATTCGTTGATGGTTAGAATCATAAACTGGGCAAAGTCGCCTTCTTCCCTTAGTAAATGAATTGGCATGCCATACCAACCATTAATTGATACTGTTTTATTTGATACTCCACTCATTGTATTAGATGGAAAAATCCCTTTACAGAAGCTAGCCTACTTGCTCGGTAAAGAGGATCTGGAATAGTTATAACGGTTGGAGAGGCAAATTGAGGGTTTTATTTATATGTGTACTGAAAATATACCAATTTTTTCAATCAAAAAACCCCGATGCGGCCGGCCGGTATATATGGTAACTAACATGAAATAATGCACCAGAGTAGTTGATGAAATGTTTCTGAAGAATAAGGCGATAAACGATAGGCAACTGTGTAGATTTAAATATTTGGCCAATCTCTATGTACTTTCTCTTTTTTTCCAGTGTCAAATACTTGTAGAAACAGTCTAATTCATTAAGAAAGTATATAAAATCTCTCTATATTATAC tpg|BK006938.2|:1050818-1053153 7X171= 518=7X 
 tpg|BK006941.2| 886850 + tpg|BK006941.2| 886868 - INS GAACATATAGTTTTATCCTTAGAAGAACTATCAATTAGATGTAGTAGCTCATCACTGAATTTTCTTTCACGTATATCATAAAGGTTCATACCACAGGCATCTGCCTCCTCTAATTCAACAAGATGGCCCACTAAGATAGAAGTCAAAAAATTAGACACTAAAGAAATGGTCTTTGTTTTTTCGTAAGCTTCTGGTTCTAATTGTGCAATTTTCAGAATTTGAGGACCAGTAAATCTAAAATGGGCTCTGGACCCTGTTAATTGAGCCATTTTTTCAGGCCCACCTATGCACTCTTCAAACTC tpg|BK006941.2|:886232-887486 7X350= 151=7X 
 tpg|BK006941.2| 984239 + tpg|BK006941.2| 984028 - INS TGTAGATTACCTCCACTTTAATCGGATGTCTTTTTTTACGTCCAAGAGTATTCAATGTCATCAAGATAGAAGCAAATTTTTCTAACACTAAATGTTATATTGCATCTGTATCAGTATATATGTG tpg|BK006941.2|:983766-984501 7X4=58S 57S5=7X 
 tpg|BK006941.2| 724581 + tpg|BK006941.2| 725018 - INS ACTATTTCTGTCGCAAAATTTCGTAAGATTTTATCGTAGTAAGTCTGAACTATATCCAATTTCATTGCCTTTGGATGGCCTGTATTCATAGGTATTTCTACTAAAATCAATCTCATGTATGGTTTATGTGACGTGGCTACAACTAGCATGGTACTGGGTGATAATCCTATCGTATCCTTAGTATTGGAATGAACATAATCTACTGCCATTACGTCTCGAATGTTGAAAGCGTACGTGCTAAATTCCGCATTGTTTAAGGC tpg|BK006941.2|:724047-725552 7X1=1I49=1X191= 210S7X 
 tpg|BK006938.2| 768660 + tpg|BK006938.2| 768857 - INS TTATACACCGTTACCAGCGTAGCCGAATCCCTTTTCACCGGTACATAGAGCTCTGAAGTTTTCTGCAGTCTTTGGGACTATGTCGTTGTACAACTTGAAAACGACACGGCCAATTGGTTGGCCATCAGCTTCGACATCAAAATAGACTTGGGACATGGTAGTATTAGCGGTTGAGTTTGGATTGAGTTGAGATATTAAATTCAAGACAAATCTTAATATAACCTATCTAGCGAAAAAGGAGGAACAAATGATGACGACAGTGGCAAAAGGATAGAAGGCTCAAGAGAATACGTTTATATTTATACAGGGAATCGAACAGACACTTGTCAGCGTAAGCC tpg|BK006938.2|:767970-769547 7X326= 317=7X 
 tpg|BK006941.2| 940697 + tpg|BK006941.2| 940836 - INS ACCACACAGTGGTCTGGTGTATTCGTTTCTGTATTGGTTGTTTCAAAAATTTGGAAAATATGCAATGTTTGCTTATTTGACAATACGGCCAACTTACTACCATTGGGGCTGAAACTCATCTCGTAAATATCCGCCTTGTCCACCCCTCTTCTAAATTCTTTGATTAAAGTACCGTTATGCGTACTGAAGATTCTTATAAGTGTACCCTGGACGGAACATGTTGCTACCATGGTGCCTTGACGGTTCAGTCTAACC tpg|BK006941.2|:940173-941360 14S79=41S 124S4=7X 
 tpg|BK006938.2| 1170235 + tpg|BK006938.2| 1169619 - INS TGTAAATATCCCGCTTTTAGCCATTGATGCGTCACCAAAAACATGGTTAACTGATTATGGCGTATTTGGGAAACGAGAATATTTAGAAAGGGTATGGGACTCTATAGAATGGAAAATTGTAGAGTCAAGGTTACCTCAACGTACTAAGATCCAAGCATTCAACACGTTATGAATGAAACTGGTAATGGGAATTTTTTCCTTTTGATATAAGTTGGTAGTCTCTGTAAATATATAAAGTCAAACTATTCGTAATGTGTATATAACGTGGTCTTAAATTATTTTTATTCGTATCTCTCCCTTTTATTTGCCTGGCTTTGGTGTCTCATAGCTTCTTTTCTCTCTTTTAAGCTCACTTTACTGACTTTTCCTGCCGACCTTTAGACTTTTTACTCTGCTCAGTAATTTGC tpg|BK006938.2|:1168791-1171063 7X357= 204=7X 
 tpg|BK006938.2| 860641 + tpg|BK006938.2| 860959 - INS TTGAGCCTCAAAATTCCACTTGTTGGTGCCGGGCTACTTCTATGAACACAATTTCAGCTAACCCGAATTCTTTACCGCTACAGCCTATAGCAAATTGACAATTCTTTGTCCTGCATACCTTTTATATTAATTTTTTAAACAAGATTTCATATACATAACGG tpg|BK006938.2|:860305-861295 7X5=75S 38S10=40S 
 tpg|BK006941.2| 557322 + tpg|BK006941.2| 557248 - INS GCTATTGTGCTGTGATTAAATCATATAGGAAACTTCTTCTCGAGAAAAAAGTGAGTTCACCCGCGGCGCTCTCGTAAAACCCGAGGGCCGATTCTTTCCCTCCGTGGAACAATCGGCCCCGCGGCGTCAGAGGGTATTATCTCCGCAAGTGATAGAACTCACATTTATTCTACGTTCTGCATGGTTTTGATTATCTTCTTTTGCACGATGTCACATACTTTTTCGATTACCGTCGCTTTACACAGTAACTGTTTAAAAC tpg|BK006941.2|:556716-557854 32S97=7S 124S6=7X 
 tpg|BK006938.2| 814944 + tpg|BK006938.2| 815165 - INS GAATCAGTTACAGAAAAGGTCCCATTTAGCGTAATTTCTTAGCGGAACTCATTAAAGAGCTCCGACGTGCAACGCGATAAAGGTTCGCCGACGACAACAAAACAATGGCAGGCAGTCATTAAATGAACGCCATCAAATGAAATATTCGTGGTAGCGATTACAATAAGGA tpg|BK006938.2|:814592-815517 7X4=80S 75S8=1X1=7X 
 tpg|BK006938.2| 233263 + tpg|BK006938.2| 233116 - INS CCTCCTCTATTGTTGAATCTACCGGGCTATCTAAAACATTTATAGGTTTGATTGTCATTCCTATTGTGGGTAATGCCGCAGAGCATGTCACTTCAGTCTTGGTGGCCATGAAGGATAAGATGGATCTGGCGCTAGGTGTTGCCATCGGTTCCTCCTTACAAGTTGCCTTATGTGTTACACCATTCATGGTTCTTGTGGGCTGGATGATCGATGTTCCAATGACGCTAAATTTCTCCACTTTTGAAACCGCTACTCTTTTTATTGCTGTTTTCTTATCCAATTACTTAATTCTCGATGGTGAGTCAAACTGGTTGGAGGGTGTCATGTCTCTAGC tpg|BK006938.2|:232434-233945 7X101= 144=1X16=1X162=7X 
 tpg|BK006941.2| 645103 + tpg|BK006941.2| 645725 - INS ATATATATATATATATATAATATATATGTAGTATACACACGTGGACGACCATTAACGAATGTTGTATATGCTTATGCGGAACCTTTGTACTCTCTTAAAATAACAGGGACAGATGAAGGTGGCAAAGCGCCGAATTCAGTGATCACTTTTTTAATATATTCTGGTGGTGTTAAATCGTATAAGATGTTGACAATATTTAACGAAGGTAACTCTTGCCAACCATCCAAAATATTTTGCCCTGGTTATAGCAACCGCGATATCTTCTATGGTCAACTCCAATTGTAGTTTATCAATCGTACCTAAATCAATACGCACTTGAATGA tpg|BK006941.2|:644443-646385 7X235=47S 365=7X 
 tpg|BK006941.2| 781989 + tpg|BK006941.2| 781463 - INS GTAATGGGCAATATTGATTTTTAAATTAACCGTAGAAAATACTAAGTGGAAAGATCCGATAGTGATGAGATAAGACTTTTAGTTATCTCTGTAATGGTGAGTTTTCGCACATCTTGCAATATTAAAAATATAAATCAATTCTTCAAATGTCACTTCATGGTCGGGTAACCAAATATGATCTTAAAAAAAATTAAGAAAAAAAAAAATTGAAAATTTTGAGCTAAGCTCATCTCATCTCATCGGCTGTAATCAGTAACACATCATTTATTACATCAGTTACAGGTATCAACATATATCTTCAAAAAGGGGACATTATGGTTTTGAAATCTACTTCCGCAAATGATGTTTCAGTATATCAGGTTTCTGGTACAAACGTTTCAAGATCACTTCCAGAC tpg|BK006941.2|:780659-782793 7X243= 371=7X 
 tpg|BK006938.2| 1034995 + tpg|BK006938.2| 1035162 - INS CAGATACTTATTCATAGCTTATAAATATTTACAGTGTTGTAACTCTAGTAAAAACAAAAGAGGTCATCTAGATTGCATTCTCCTTATTTTATCACTGATATCGTCTTCTTCAAGAAAGTGCAGGATCTTGGTGCACGACTTAGGATCACCAACTTTCTCAATATGAAGTACTGGTATGTCGAAGCAATATTCCTTCCACCATTTTGCGTTTCTTCGGTCAGTTATGTTG tpg|BK006938.2|:1034523-1035634 229S38= 115=7X 
 tpg|BK006941.2| 387527 + tpg|BK006941.2| 387512 - INS TTACCCCAACTTCGAAGGTCGTTGGTGATCTGGCACAATTTATGGTCTCCAATAAATTAACTTCCGATGATGTGAGACGCCTGGCTAATTCTTTGGATTTCCCTGACTCTGTTATGGATTTCTTCGAAGGCTTAATCGGCCAACCATATGGT tpg|BK006941.2|:387194-387845 7X4=72S 72S4=7X 
 tpg|BK006938.2| 1115667 + tpg|BK006938.2| 1116283 - INS ACTGCTCTTAGTTGAAGTAACCTCCAAAAGTTCAACTTCTTGCGGTTTTTCATCTTCTTCAGATTCTAGATCCACAATAAATACATCATCTTCGCAAGAGCATATGACAATTTTGGAATTATCGATGAACTTGACTAATTTTGTGGAAGTTCT tpg|BK006938.2|:1115347-1116603 7X4=72S 71S6=7X 
 tpg|BK006941.2| 345146 + tpg|BK006941.2| 344982 - INS TCTCTGCGCGTTGGCTTTTATCC tpg|BK006941.2|:344922-345206 7X4=7S 7S5=7X 
 tpg|BK006938.2| 52116 + tpg|BK006938.2| 52889 - INS CACCAGGGTTCACTTCAAGGAGGAGCTAACTCAATTCAGGAAAAATATTATGTTTGATGGGGAAAGATACAACGTCCCAATTTACAAATTTGAGGTTGACCCTGAAGATGATGATTTGGAATCCATGGAAGAGAATCAAGCCTTGGCATCCTTGCAACCATTTGCTATTATAACTTCAGATACCAGAGATAGTGAAGGTAGATACGTTAGGGAGTATCCGTGGGGGATAATATCAATCGACGACGACAAAATTTCGGATTTGAAAGTTTTAAAAAACGTCCTGTTTGGTTCTCACTTACAAGAATTCAAAGACACCACGCAAAATTTGCTTTACGAGAATTACCGTTCCGAAAAACTATCGTCCGTGGCCAACGCTGAAGAAATTGGTCCTAATTCTACAAAGAGACAGTCAAATGCTCCAAGTTTAAGCAACTTTGCCTCTTTGATAAGCACTGGTCAATTCAATTC tpg|BK006938.2|:51166-53839 7X149= 1S44=1X408=7X 
 tpg|BK006938.2| 1360888 + tpg|BK006938.2| 1361216 - INS GTAAAGTACCGGGAATGCTTTACAATGAATCAGCTATTGGCGGATATTGACCAACCAACACTAAAATTTTATATCCTGCTCCGATTTTTGTCTTGGCCGTGAAATCCATTATGCACATTTTTTACTAACGTTTATCAATAAGTTCGGTTTCCCGTCTAAATTTTTT tpg|BK006938.2|:1360542-1361562 7X4=79S 77S6=7X 
 tpg|BK006941.2| 774842 + tpg|BK006941.2| 774708 - INS GTCAACATTCGCTCGAAAAAACAACCCATATTCCATTTGATTCTACGCAGCTGGTAGAAACTTTTACAGGTTTGATAAAATTATTACAATCGTTAGCGGTTACGCAAGGAATAGGAAATAAAGAAACGGTAAATAATAAGAAAAACACAGCAGATCTAAGCCTATTGCACACAGTATATT tpg|BK006941.2|:774334-775216 7X373= 158=7X 
 tpg|BK006938.2| 1377281 + tpg|BK006938.2| 1377276 - INS CTCCAGAGATGAATACATTTTTATTTATACTAAGTGAAGGTATCATAGATCAGCACTCTTTGGAAAAGGTTTATAACATTATTTCCAGCAGGGCAATGGGGCACGCAAAAACCACGACCGTTAGACAGTTACCATCAGATTGTACCCCGCTAACAGTGGCTAATCAAACTATCGAAATTTTGCAAAGTCTAATTG tpg|BK006938.2|:1376872-1377685 7X5=194S 98=7X 
 tpg|BK006941.2| 1082414 + tpg|BK006941.2| 1082503 - INS GATAGAAAAAGGGCAACAATGTTGAGCTATTTTAGGCACAGAAACTTTACTATTCGAAAAGGGCATCCATTTCATTTCCGATTTTCTATCTAGCTCACTCGATAATCGTAATAGTACTTTTATAAAACTTTAGTGCGGGTACTGTGAGAGTG tpg|BK006941.2|:1082096-1082821 7X4=72S 71S5=7X 
 tpg|BK006941.2| 596926 + tpg|BK006941.2| 597187 - INS CTTGTCTGATGAGAACCTACACTATTATGGTGAAAACACACTATACTTACTGTCTTTCCAAGGTGTCAACGGGACTTTGGGTGGTAACTCTGTACGTGTTTCTTTAACCACTGGACCTGTCCACGATTTCACTTGGTCGCCAACTTCAAGGC tpg|BK006941.2|:596608-597505 29S30=24S 73S3=7X 
 tpg|BK006941.2| 177459 + tpg|BK006941.2| 177373 - INS GTTGGAAAACCATTGTCTCATTGTACTCCAGTGAACTAGTAAATGGTAAAGACAATAACGTGGGGAAACCCGCCAGCATTTCGGCACCGAGTTTAGCATTAGGTAATAAACCATAC tpg|BK006941.2|:177127-177705 7X4=54S 53S5=7X 
 tpg|BK006938.2| 664851 + tpg|BK006938.2| 665308 - INS ATATATCATTCCCGAGATATATAGCACCATTAGTATTGGTGCCTTGAAAAGCACTATTAGCAGCGGCTCTAGTTGTGGTGTAAGCAATCGCAATAAAAGTAAATAAAGAGCCCAAAATGATACTAAACTTACGGGTTCCACTAGATCTAACCAACGGATTACACATTTTGTCATCCGGTTCGGAAGACATGGCACTCATTGTCAAATAAGTACAGTAAACAGAAACCATACTACTTTGGGCCAGCCCACTTTTAGGGTTGGCCTCTTGGATCTTAGGATTCACCGATAAGACAAGCGTTATAAC tpg|BK006938.2|:664229-665930 9S170=56S 70S6=7X 
 tpg|BK006941.2| 522883 + tpg|BK006941.2| 523416 - INS TTAGCTGATACTAAACGAAGATTAGAAAAAGAGCAAAAAAAAACAAAAAAAGAACCACCGAAACATTAAAAGTGGGAATAATGTCGCATCAAATGGCGCCATGGATACCCATGTTTATTCAATCGTGCAAAAATAACACTGAACCGTTTGTATCATTTCAATTTGCTACTGTTGAC tpg|BK006941.2|:522517-523782 7X76=56S 1=246S 
 tpg|BK006941.2| 662759 + tpg|BK006941.2| 662295 - INS AAGGATGTACTAACACTTTGTGGTAGAACATTATATTTTTCATAGAAATTTTACAAAGGATCTCCTTCATATACCATGGCTACAAGTGTTAAAAGAAAAGCATCTGAGACTTCTGACCAGAATATTGTTAAAGTGCAAAAGAAACATTCCACACAGGACAGCACAACTGACAACGGATCCAAAGAAAATGATCACAGTAGTCAAGCCATCAACGAGCGTACCGTGCCCGAGCAAGAAAACGACGAAAGCGATACTTCACCTGAAAGTAACGAGGTCGCTACTAACACTGCTGCGACTCGCCACAATGGAAAGGTTACTGCAACAGAGTCCTATGATA tpg|BK006941.2|:661607-663447 7X4=250S 3S7=1X14=1X301=7X 
 tpg|BK006938.2| 1395947 + tpg|BK006938.2| 1396648 - INS CATTCAATGCCGTGAAGTCTTCGACAATAAATAACAATGAAAATTGGGTCGATTGCTTTTTCAGAGCAAGACAACTACTAGAAGAAAAGCAAATTCTTGATAAAATCAGTAACGTTTCCTTTGATAGTAAGGCATCGAGTGAACCATCATCACCTCCGCCTATTTCAAGAAAAGAGCGGCCTCTGAGTATAGGAAATAATGTAACAACACTCAGCTATAC tpg|BK006938.2|:1395493-1397102 7X82=28S 2S1=188S 
 tpg|BK006941.2| 514132 + tpg|BK006941.2| 513658 - INS GTTAAATCCAAACCAATACGTAAATGCCGCCAAAAAGGCATGTAATGAACTAAAGAAGAGTGGTAATGGAATAAGAGCAGTTTTTGCCGATCAGTTCGAAAACGAAGCCAACTGGAAAGTACATTACCAGACCACAGGCCCAGAAATTGCCCATCAAACTAAGGG tpg|BK006941.2|:513314-514476 7X5=161S 83=7X 
 tpg|BK006941.2| 690355 + tpg|BK006941.2| 690476 - INS CAGGAGCAAAGGATTCCGGGAGATTGTTTTTAACACCTCATTTTCTGGTATTTCGAGATGCATTTGATCATTCATCGTGCGGACTAATACTGAATATTTCTACCATTAAACGTGTAGAGAGGTCGCCATCCGAATCATATGAATTTGCTCTTCTAGTAACTTTGTACACAGGAGCAAAGGTTCTGATTCAATTTATCGGTATACGTTATAGATC tpg|BK006941.2|:689913-690918 7X165= 55=1X132=7X 
 tpg|BK006941.2| 1027813 + tpg|BK006941.2| 1027763 - INS CTATCAGGGAAAAAAGATTTCTTCGCGAAAGAACTAAGCCGGTAAATTACAAATTACCACCACCACTAACTGCTAGCAACGCAGAAGAATTTATAGATAAGAATAACAATGCACTTTCTTTTCATAACCCATCACCTGCACGGCGTGGTCGCGGTGGTTGGAATGCTAGTCAAAATTCTGGTCCCACAAGAAGGCTTTTTCCCACTGGTGGACCTTTTGGTGGCAATGACGTAACTACAAT tpg|BK006941.2|:1027267-1028309 7X162=18S 4S1=254S 
 tpg|BK006938.2| 893650 + tpg|BK006938.2| 893907 - INS AAGGAACATGCGGAACATGCTAGAATGATTGCCGAAAGGGCGGGCCCTAGTCAATGGCATCATGCGGGAACGTGCAGTAAAGCTCAATGTAACTTGATGCCTATCGGCGTTGTTCGAGCTAAGGACGATGTGATAGACTGAGGAAGGGTGAACGTCGATAGTTAGCCGTTGTGAACTAAATAAAAGTGATATTTTTTCGTTGTTCTTTTCTTGGT tpg|BK006938.2|:893206-894351 7X80=27S 3S1=445S 
 tpg|BK006941.2| 237898 + tpg|BK006941.2| 237216 - INS GTTTAATACATGTCGATAATTGCATTTGCAGTAAATACCAGAAAAAAAGACCGTAAAACTTTGGAAAATGTGATGAAAAGTAAATGATACTGCTTTTTGCCTACCAAGTTTAATATTAGGGAAATGCTGGGAATTACCCAAATAAGTCCACTGCTGGGTCTTTGCAAACATGCCAGAAATGCAAAAATAAGCGACTTAGTAAAAGATGACTCTTTTATCATTTGTCCGCCTGTCCAGTCCCAGTAGTAGAGGGCAATAGAAGTTAAAATCATTTCAAAAGAGTTGATGAACGTTCTTGTAATAAAAAAGCAATTAAAAAAATTAGTTAAACTTAAAAGC tpg|BK006941.2|:236524-238590 21S15= 170=7X 
 tpg|BK006941.2| 913639 + tpg|BK006941.2| 914364 - INS GCCCACACCATGTGGCAAAAAAGTCAACAACGACTAACTTGTCGCCAGATGCTAAAGCACTGTCGTATTCAGAAGCGGATTTTAATTGAGTGAACATTATTGATGTGTTATTTAAAGATATCGTAGACTCTCGTGTATGTGTGCGTGTATAATTCTTGCTAGACAACAAATAAAAACTGGTCCTCGTTATTCTCTTGTCAGCTTTTCATCCCCCGAATGGCTTTCTTATATACTGATATCCCTCTTT tpg|BK006941.2|:913131-914872 7X2=181S 124=7X 
 tpg|BK006938.2| 290510 + tpg|BK006938.2| 291247 - INS AGAGTATTTCTTTGCCAAATCCAGAGAAGGTTTCTTATAAGAAAATGAGCTTTTGGCAGAAGTTTGTTGCTATCCACAAGTTCATGTTCTACCTTAACAATTATATGGATACTAGTCATGCCTACTCATCTGAACCAAAGACTTGGCCTCTTATGTTGCGTGGTATTGATTTTTGGAATGAAAATGGCAGAGAGGTGTACTTTTTAGGTAACGCTGTTTTGTGG tpg|BK006938.2|:290048-291709 7X246= 112=7X 
 tpg|BK006938.2| 214424 + tpg|BK006938.2| 214582 - INS GGGTGGTGTCAGATCGAAATGTACCGCCATATGCGCTGCCGCAAATTGGCTAGTTAATTTCACCTGTGCCCTGATTACACCTTACATTGTTGATGTCGGATCACACACTTCTTCAATGGGGCCCAAAATATTCTTCATTTGGGGCGGCTTAAATGTCGTGGCCGTTATCGTTGTTTATTTCGCTGTTTATGAAACGAGGGGATTGACTTTGGAAGAGATTGACGAGTTACTTAGAAAGGCCCCAAATAGCGTCATTTCTAGCAAATGGAACAAAAAAATAAGGAAAAGGTGCTTAGCCTTTCCCATTTCACAACAAATAGAGATGAAAACTAATATCAAGAACGCTGGAAAGTTGGACAACAACAACAGTCCAATTGTACAGGATGACAGCCACAACATAATCGATGTGGATG tpg|BK006938.2|:213584-215422 7X177= 23=1X183=7X 
 tpg|BK006941.2| 525196 + tpg|BK006941.2| 524718 - INS ATATTTGTATATGCTTTGTATTCGCGCTATCTCGATTTCTACCTATATAGTTAATCTCTGTACAAAAACAATCTTTCCAACTATCCATTAATCATAGTATATTATCAGCGTCGGCGATTTTACCACGCTTGACAAAAGCCGCGGGCGGGATTCCTGTGGGTAGTGGCACCGGCAGTTAATCTAATCAAAGGCGCTTGAAGGAAGAGATAGATAATAGAACAAAGCAATCGCCGCTTTGGACGGCAAATATGTTTATCCATTGGTGCGGTGATTGGATATGATTTGTCTCCAGTAGTATAAGCA tpg|BK006941.2|:524098-525816 7X4=33S 285=7X 
 tpg|BK006941.2| 220755 + tpg|BK006941.2| 220791 - INS GTACTATATGATACTTCTGCATGAAAGAAAATTATTGAATGATTTAGCGTTGGAAAACGGCGAAATAACCAAGACAGAAAATGAGAAATTTATCAGTTATCACGATAAGTACTTGTGTATGCTGAAAACATGCGTATTCTGAGCCATCTCTCCTGATATATAAGAC tpg|BK006941.2|:220409-221137 7X9=146S 28=1X117=7X 
 tpg|BK006941.2| 934857 + tpg|BK006941.2| 935208 - INS AAAGGTTGGGCGTTCAAACATAACAATAGAGATGTCGAAGTTAATGGTCTACAGATTGCATTAGAC tpg|BK006941.2|:934711-935354 7X10=138S 33=7X 
 tpg|BK006941.2| 960671 + tpg|BK006941.2| 960683 - INS GTACTTGCGCAATAAATAAAGAGTTGATACACCAAAACGAAGTTCCATTGGTGTTACTATCGTCTGGTGTTGGTGTTACAC tpg|BK006941.2|:960495-960859 7X3=113S 41=7X 
 tpg|BK006941.2| 179364 + tpg|BK006941.2| 179387 - INS ATGACGAACATGTTCAAGCGATTTTTTTTCACTATTTCTTCTACCAAATGTCACTTCTTCTCTCAATAACGCAAAATGTGGCCCATGAGTAGACAAACCCAGCATAATCAAATCTGCGTCAAGACCGTAAATACAATGTCTCGTATTCTGGTTGAAATCCTTTTGGGATTTTAAATGCCTTATAAAGTTCATGATCTTGTGTTCACCTTCACCTGGAACTTCATGGCCAGAAAATATGATTTGCACTTCCCTCCATTTGGAATCGTTAGAAATCTTGTCGTGAATAAAATATTGTAAGTTTTTGGTCAATTTGGCCATAAAC tpg|BK006941.2|:178706-180045 7X171= 302=7X 
 tpg|BK006938.2| 1068160 + tpg|BK006938.2| 1068226 - INS CTTTATGCCAGGGTAAGTGAACAATACATATAAAGGATATTTAATGCTAACTAGCCCGATATATACATCTATCTATCACTAGGCATTCGAGTAGTGAATAAGAACCACTACTTGAAACACTAGATTTGTAACAATAACGCATGTATCATCGTACATTTTCG tpg|BK006938.2|:1067824-1068562 7X6=74S 71S8=1X1=7X 
 tpg|BK006941.2| 646967 + tpg|BK006941.2| 647130 - INS GTTCTACCTAATGTTGCAACAAGAATATTTGCTAGTCCAGTATTATTTTTTCTATTTAATACCTTTTTCCAAGCAACCTGCAGTTTCCTCTGAGCAATTTCTGCATCTTTATAGTCTTTCAACCTATTTCGATGCAAAGCACACATGATATTAGTATTAAAAAAATGCTCGATATCAAAT tpg|BK006941.2|:646593-647504 7X1=1I73=15S 17S1=279S 
 tpg|BK006941.2| 293239 + tpg|BK006941.2| 293139 - INS TCGCTATAGGGTCTCTGGTGCTAACATCAAATTTTCAATTTGGCCTGCAAACCGGTTGGGTTTCCATGATGTCCCTGCCATCGGCATTGTTAGCTTGTGCTTTCTTTAAAAATATCTGGCCATTAATATTTCCGAACGACAGGCCTTTCAGTGACGTTGAAAATGTATACGTACAAAGTATGGC tpg|BK006941.2|:292757-293621 7X65=27S 9S1=104S 
 tpg|BK006941.2| 882688 + tpg|BK006941.2| 882859 - INS GGTGAATGCAATGATACCGTATTCGTTGTCGTACCAGGAGACCAACTTGACGAACTTTGGAGACAATTGGATACCAGCGGAAGCATCGAAGATGGAAGAGTGAGAGTCACCCAAGAAGTCAGAGGAGACAACAGCGTCTTCGGTGTAACCCAAAACACCCTTCAACTTACCTTCAGCGGCAGCCTTAACAACCTTCTTGATTTCATCGTAGG tpg|BK006941.2|:882250-883297 7X4=76S 2S197=7X 
 tpg|BK006941.2| 373608 + tpg|BK006941.2| 373603 - INS TTGTTCCTCTATACTCTTCTCTCCATTAACTACAAACACGAATAATGAATTTGAAGGAGAGTCAGATGA tpg|BK006941.2|:373451-373760 7X3=31S 31S4=7X 
 tpg|BK006938.2| 465337 + tpg|BK006938.2| 465808 - INS ACCCATGACTAATAGCGGACGTACCCGCAGAGACATAAAAAAAGAAAAACTATATCGAAGACCGAAAGCAGTAAAAAAGTGGATAGAATAACACAGCTACCAAAATACGGAAAGAGAATTCAATGAGCAATATCAAAAGCACGCAAGATAGCTCTCATAATGCTGTCGCTAGAAGCTCAAGCGCTTCTTTTGCAGCTTCAGAAGAATCATTTACGGGCATAACCCATGACAAAGATGAGCAGAGCGATACCCCGGCGGATAAACTAACAAAAATGCTGACAGGACCTGCAAGAGACACTGCGAGCCAGATTAGTGCCACTGTGTCTGAAATGGCGCCAGATGTCGTATCTAAAGTGGAGTCATTTGCAGATGCACTATCCCGTCATACAA tpg|BK006938.2|:464543-466602 7X201= 97=1X280=7X 
 tpg|BK006941.2| 716560 + tpg|BK006941.2| 716336 - INS GTGGAGAAGGCCATAGAAGAGACAAAGCTTCATGGATTGCAAGAATTAGAATTTTGGGACGAAGAAATTCCCATCAAAAAGTACCCACAATTGTTTCAGTTATTAACAGAGCTTGAAAATGAATCTAAAGTTTTCTCAGAAAACGGTTCCATCAGTGCTGTTCGTCCCCCCAAAGGATATACAGCCGAGCAGGTAATTTGGGATAACAATACCAAAT tpg|BK006941.2|:715888-717008 12S198= 9S5=7X 
 tpg|BK006938.2| 454102 + tpg|BK006938.2| 454660 - INS GTGCTAACCACATCATTGCTCCAGAATACACTTTGAAGCCTAACGTTGGTTCTGATAGATCTTGGGTGTATGCTTGTACAGCAGATATTGCAGAAGGTGAAGCAGAAGCCTTCACTTTTGCTATCAGATTTGGCAGTAAGGAAAATGCTGATAAATTT tpg|BK006938.2|:453772-454990 7X5=74S 72S7=7X 
 tpg|BK006941.2| 314397 + tpg|BK006941.2| 315017 - INS AGGTTCACTTGCTAAGGATTTGATTGTTCCAAGGAGGCCTGAATGGAACGAGGGCATGTCCAAGTTTCAGCTTGATAGGCAAGAAAAGGAAGCGTTTTTAGAATGGAGAAGAAAATTGGCACATTTACAAGAAAGCAATGAAGACTTGTTGTTAACACCGTTTGAAAGAAATATCGAAGTTTGGAAACAGTTATGGAGAGTTGTTGAAAGATCAGATTTAGTTGTTCAAATTGTAGATGCGAGGAATCCGTTGCTGTTTAGATCTGTCGAT tpg|BK006941.2|:313841-315573 7X161= 136=7X 
 tpg|BK006941.2| 1015070 + tpg|BK006941.2| 1015368 - INS TTTCTGTCATGGTTACCGTTCTAACCAATGCTTCAATAAATTTAGTATTTTTCATCTGCAATGGTGAAGCTAACTGATATAGCGCATTGCAACACGATAAAATCACTGTAGGGTTGGAACTATAAATTAAGCAATTCAAACTCTGTAGAAATAAATCTAAATCAGGGTCATTTACCACCTCGTAAGATGGGTATTCAATCTCGTTGTATTTATCTGGTAAAGGACAACTCCTTGGGGAACCTTCTGATGATTTATCGACCACAGTTGGTTTTGGTAAATACTGCTT tpg|BK006941.2|:1014484-1015954 7X258=10S 4S1=161S 
 tpg|BK006941.2| 928539 + tpg|BK006941.2| 928586 - INS TTTGGGCATAGGTGCCTCTATATCGTATGC tpg|BK006941.2|:928465-928660 7X4=11S 11S4=7X 
 tpg|BK006941.2| 659197 + tpg|BK006941.2| 659057 - INS AAGTGAGACTCACTGAAAAAGAGCTTGAATTAGAAGAGGAATACTTGAAAAAGAAAGATCTACACTTGAAAAATCAATTAGAGTTCAGTAAGTTAGAAGAAAGCTTATCGAAAGACCTGAAAAACTCAGAAGGGAGGTTCCAAAAGGTCAATCAAGAATTAGTTCAACTAGGCTCTAAACTGGACAAATTGAACGCGAGAAACGAGAAGTTACAAAAGGAGGTCGATCAGAACGCAGAAGAGATAGAAAAGTTCAGTACTCAATTTTTGAGTAAAAGAGAAAAGGATAGATTTAGAAGAAAGGAGTACAGGATACGCGAAGCCAATAAATTTGAATTGACTATAAAGG tpg|BK006941.2|:658347-659907 7X1=1X9= 327=7X 
 tpg|BK006938.2| 903678 + tpg|BK006938.2| 903758 - INS CATCGTATCTAACGCTAACAAGGCCGTATATTTATTTAGACCTTATTTGGATGGGGAGCTGCCAACATTTTCTCCAATAAATCAATCTTCCTTTGATAGTCTTCAATAATTCTGTTTTTTTCGTCTATTTCTTTGTGTATTTGATAAGCATTTTCATCGTTTGTATCTGGATTCCCAAGTGTTCTACTTGCACTATTTCTTCTGGTGGAAACATTGCTGACACTTCCCCTTGAGGTTTCGTCGATAT tpg|BK006938.2|:903170-904266 7X222= 124=7X 
 tpg|BK006941.2| 811406 + tpg|BK006941.2| 810715 - INS ACATTATACCACGAAAATCCAAGATTTGTAAAATATGAGCCGCGTATTTCTGCAATGGTAGAAACGATAATGTACCTATCGTACAACGATACATTATTTTAGTGCATTATAAGCCGCTTGATTCATGTTGATAATTAGCGGCTAAATTGTAGTAGTCATTCAAAATAATCGTACACCTTCATATAGTTATGAAAGGGGTATAAA tpg|BK006941.2|:810293-811828 7X5=4S 102=7X 
 tpg|BK006941.2| 432597 + tpg|BK006941.2| 432612 - INS GTTTCAGCAATGGGCGTGTTGGAATTTTCTTTCGGAGCAATAGCAATAGGAATTAAAGGCGATAGGTGTTGCTGTGGTAATGGCGGTGAAAAATTTGCCGTATTTAAATCTGGTATACTGGTAGCACTAGAACTAGCACTATTTATTGGAGAGCCCACAACCTTCTTCTTTCTGCCTCTTTTACCTCGAGGGTGGGAGTTTGTATGAATTCTTCTGTGTCTCGTCAGTTCATCGCTTCTACTGAACCTTTTCACACATCCGGGGAAGTCACACGCG tpg|BK006941.2|:432031-433178 7X5=248S 4S255=7X 
 tpg|BK006941.2| 246013 + tpg|BK006941.2| 246039 - INS ACTTCCAATCTGTTGTCGTGGTTGCCATGCAACATGTTCATCGAGTTCCGCCTATTGCAGCCGCCTGGGCGGAAAACTTGGTTTGGTCAATGGGGTTAATTAGAATCTCATTCATGCAAAGGATTTTCCGGTGGTATGTGCAATCCACTGGTGGTACGCCTAGCTTATATC tpg|BK006941.2|:245657-246395 7X46=39S 2S1=28S 
 tpg|BK006941.2| 958187 + tpg|BK006941.2| 958867 - INS TTCGTATAATTGCCAAGACATAATCTAATTGAGAAGGTCAGACGGCAAAACAAATGACCGAAATCTTCGTTTATTGGTTCGCCTGCGTTGCCAACTGGTACATTTTCCCAGAGTACCAGCAAAGGAAGGCATCCTTGATGCCTACTCTGATAC tpg|BK006941.2|:957867-959187 7X5=71S 73S4=7X 
 tpg|BK006941.2| 861677 + tpg|BK006941.2| 861047 - INS GGGTAAGCTAGATCATAAATAATACTTTCGGAGTCCAATCCCTCCATTCGTACATCAGATATGGTCCTTAGGGCGAAGAGCATCTGCTCACTTACTTTAAGAACATCCCCAATTTTGGACGCTTTAGCATACAATTTGGTAACCTGTTCTGCATCAGAAAGACCCTGAAGAAAATCTCTTAGAAACTGTCGAGAGAACGTTGTTAACGCCTCTGTAACAGTCTGACGAAGTGAAACTGGAGAAAATAAAGCGCTTCGAACAATATATTGGAAGAGTTGATTTTGGTTCCAAACAGTATCGGGC tpg|BK006941.2|:860427-862297 7X6=4S 39=1X112=7X 
 tpg|BK006941.2| 670662 + tpg|BK006941.2| 670827 - INS TCCTAGTGTATTTAACCACAGCGAAGGGACCTTTAAGTGTTCCTAAGGGTGATATGGATATCTCAGGCCATTGCCTCATTATTCCCATTGAACATATTCCGAAATTAGATCCAAGCAAGAACGCAGAGTTGACACAGAGTATTTTGGCTTATGAAGCTAGTCT tpg|BK006941.2|:670322-671167 7X4=77S 78S4=7X 
 tpg|BK006941.2| 326767 + tpg|BK006941.2| 327177 - INS AAAGCAATGTTCATCTAAAAACACAAGAAAACCCTCAAAAAGAGTTATTGTGTGCAATAACACTAAATGGACCACAGATACATTTTTGAAAATGATACAATCCGTTTTTGCTTATAAGTACACTGAAATAAAACCTACCTGAGCTGGCGGCGCTACAAACACTCAATGTTTCTAACATATGGAACAAAGAGAAGACAGCAAATTACCTTGCTATAAC tpg|BK006941.2|:326319-327625 7X123=39S 1=21S 
 tpg|BK006941.2| 56986 + tpg|BK006941.2| 57230 - INS GCGTTGAAGACCATAGATTCACAGATTGTGAAGCCGACGATTGATGGGATGAGACG tpg|BK006941.2|:56860-57356 7X4=108S 7=1X20=7X 
 tpg|BK006941.2| 558163 + tpg|BK006941.2| 558344 - INS ACGCACCGAACGATACGGGGCGTGGCTGTTTTATTATATTCTTGATCACGTTATTGAATATTTCGTTCATCAATTGGCCAAAGGCTACAATGCAGGCTTCTAACTCTCTTGTGATGATAAACCACGACAAATAAAAAGCTAGCACTAGGATGGGCATCAGCGAGAAATATGCACTAAGGAATGATAGAAAGTCATGCGAATCATAGAGAATGTATGTG tpg|BK006941.2|:557713-558794 7X200=4S 6S1=248S 
 tpg|BK006941.2| 89348 + tpg|BK006941.2| 89218 - INS AATCTAGAAACATATTTTCCTAAAATGAAAATCGGAAGCTAACAAAATTTTTGAAAAACGAAATAAAGAAGAAAGATTATTATTATTACTTTTTTTATTAGTACTCCATATGGACCTCTTAGGTG tpg|BK006941.2|:88954-89612 7X109= 179S1=4X3S 
 tpg|BK006941.2| 719075 + tpg|BK006941.2| 719788 - INS GTATTATGAGTGGTCAATGGGCCCGTTACGAAGAACAGAAATTCAATGTTCTCAGGACGTGCTGAAAGGAAACCCACAGAAAGCAGACATTCTGTTGCAAAGAAAACTGAAAAAAAAATAAATACAAGGCCCCCCTTCAGATGACTACGCCCAACCCAACCAAAGAATTATCCTCCTCACAAAATATATCGCT tpg|BK006941.2|:718675-720188 7X227= 97=7X 
 tpg|BK006938.2| 1479162 + tpg|BK006938.2| 1479737 - INS ATATGGCAATCTCCCAACAAGCACCCGCTCATATAATACCATGCAAGTGACCACAAGATTTATATCTGCGATAGTCTCGTTTTGCCTGTTTGCTTCTTTCACGTTGGCTGAAAACAGCGCAAGAGCTACGCCGGGATCAGATTTACTCGTTCTAACAGAGAAGAAATTTAAATCATTCAT tpg|BK006938.2|:1478788-1480111 7X6=84S 84S6=7X 
 tpg|BK006941.2| 806256 + tpg|BK006941.2| 806962 - INS AAAGATAAGTTACCAACGAAAATAGTAGCTGGTTCTTCGGTTTCTTCATTTTTTTGCTTCTTGTTGGAAGACTCTTCGTCTTCTTCTTCTTCGGCGTCCTCAGATTTACGTTTCTTATCGTTAGACTCTTCCTTTTCGCTTTCGCTATCAGAAGATGAAGATGAGGATGAATCAGAGCTAGAA tpg|BK006941.2|:805876-807342 7X12=156S 161=7X 
 tpg|BK006938.2| 27362 + tpg|BK006938.2| 27866 - INS TGGCAGGATATCATTTATTCATTCTTTCGTTGTGGAATTCCTTCTGCAAGTCTTCTATTCTTTGAAGTTTAGCATCATTCATGCTATTAAGTTCTTCTAGTTCTTGAATCCTGTCATCCTTCTCTTCTAGTTTTTGTCTTAGTGCTTTGATCTCTTCATTTTGGGACTGGAGCTCATCTAATACCTTGGGTAAACTATTTTCTTTAGAAATACTTCCTCCATATGATGAAGAAGATAGCCTAATTTCTCCTAATTTCATATATTCGGACTGTTCTTCATCTGGAGTTTTAGATGAGCGAAATACGTTCTCTAGATGCGCAACCTCTATATTCT tpg|BK006938.2|:26682-28546 7X151= 1S312=7X 
 tpg|BK006941.2| 727951 + tpg|BK006941.2| 728678 - INS GGCTTAGACCAAGCAAATGATGGTTGTGTGGATACCGTGTTTCCAAGTCCGGGCGCAGTGTTTGTTTGAGGCTGCTGGGATTGGCCAAAAAGGCCACCTCCCCCAAGGGTATTGTTATTCTGGGTGCCGCTTCCAAACAGGCCACCATTAGTTGTTGATC tpg|BK006941.2|:727617-729012 7X93=27S 1=166S 
 tpg|BK006938.2| 929785 + tpg|BK006938.2| 930002 - INS CTTGTGCTTAGGCAGTCTTTCTTATGTGGGCTTGGAAGACTGGTAGCTGTTTCAAAGCTTCATCGATATGAGGCTTAATAAAGCCGGCGATATTTGGACATTCTTTAGGACCATACTTGGTGATTAAACCTTGTCCCAAAAAGAGCTTGGATACGAATTCAATAGATCCTGTTGTGAATAAGATAGTGTAGGCAACCTTCAAAAAGAAAGTGATCAAGTTAACTTTTTTCAAAATTAACAAGGCTAACAGAGACCCACCGAAATATTTACCGGTTTGAACAGGGTTCCTCCATAATAGCAAATCGCAATTACAGCTTTTTTGTTGTTGTTGTTGTTGGGCTTGGCTATGTTGAGCTGAGGCGGACATATTTGCGTGTGTGAATATATATTATATATATATACG tpg|BK006938.2|:928965-930822 7X207=1X20= 378=7X 
 tpg|BK006941.2| 701105 + tpg|BK006941.2| 700537 - INS CCGTAATATGGCATCGTATTTTAAAGGAGTTAGATCGGTTTCAAAAGGTCATGCTCCGGAGTAATTGACTTGATTTTGCAAAGCTTCACTTAAATGGCGTATCTTCCTTTTATAAATTGCGTTTGCTTTATTCCCTTACCCAACAGATGAATTGGTACTCTGGCCGAGTGGTCTAAGGCGTCAGGTCGAGGTCCTGATCTCTTCGGAGGCGCGGGTTCAAACCCCGCGGGTATCAATATTTTTTTGAATCTACGCACTTCAATAA tpg|BK006941.2|:699993-701649 7X6=97S 249=7X 
 tpg|BK006941.2| 248978 + tpg|BK006941.2| 249182 - INS CTCCTAAATCCTTTTGAAAGGGTAGAATATGATTCCAAATTGGCTTTCCTCCTTTACAAAAGGTCACTTGAAGAAAATTATTGATTTGCAAGGGCGCTACCTGGTATTCATATTGTTTTTCAATTACAAAGCCTGTGTACAAAGTACTTTGTTTTTTGTATTGTTCGTACTCCTGCTTCAAGTTCTGTAACTTGTCACCTTTAAGAACATTTAAGAAGAACTCTGTCTGGAAATTTTGGTCTTCGAACTTACACACATCATGTCCAGGAAATGAACTTTTTCCTTGAACGAAAGTGCTCTTAAATAAGG tpg|BK006941.2|:248346-249814 7X1=1X9= 155=7X 
 tpg|BK006941.2| 668622 + tpg|BK006941.2| 668954 - INS GCTATACACATC tpg|BK006941.2|:668584-668992 7X5=1S 1S5=7X 
 tpg|BK006941.2| 1043617 + tpg|BK006941.2| 1043881 - INS CTGCTTTACCATATCGCCTTATACTCCTGTTGTACTTCTTTTTCTCTCTGTGTTTAAAATGCTATTTATTCTCTTAAAAGCACATTTGAAAACCATCGCCGCGAAATGAAATTATCGACTAGTTTATTAATGAACAAGGCGATAAAACCTAATGTTGGAAAGAA tpg|BK006941.2|:1043275-1044223 7X5=77S 75S7=7X 
 tpg|BK006941.2| 760505 + tpg|BK006941.2| 760236 - INS CTTCTGATACTATGCAGCATGAGGGCAGGAAGAACTCTGACATAGAGAAGAAGCTAAACGCTAAGCCAGCTTCTGAACTGAATCTGAAATTGTTAAACCTGTTTCCCTCAAAGCCTGCAAACAAAGACGATAGTTCCCCTATTAACACGTTGCGTAGT tpg|BK006941.2|:759906-760835 7X4=75S 75S4=7X 
 tpg|BK006938.2| 1434756 + tpg|BK006938.2| 1434577 - INS ACCTTGTGGAGAAGCCTGTAGTTCAGACCCGCTCTGAGAATTGCTGCCATCTACGAAAGGACGAGGATACTCTTGCGTTTGTGTATGTTCCGCAGATGTCGGTACCAAGGGCTTGGACAGCAGGGCGTGGTCTGCCTCTGTCAAAGACCTATTTCCCATATTAATGATATAGTAGCAGTATTCAAGCAAGTACACGTGCGCAAGTTGTACCAGATAGTGACTGTCCAGCG tpg|BK006938.2|:1434103-1435230 7X5=231S 115=7X 
 tpg|BK006941.2| 1050194 + tpg|BK006941.2| 1050357 - INS ATGAGAAGATCCTATTGCAGCAGGGTGTCGCGCGAAAAGCGGTGCCTACAAATTACAAAACCCTCTGGGAAATGACCGTGCAGGGTCGTTTGTGGATGCATCTCGATTAGGCCGGGCTAGGCATCTTGATTCTTTCCCAAAATGGAGTTAACGAGCTCGATTGGGCGTTAATTGATGGATTTGGTTACAC tpg|BK006941.2|:1049800-1050751 197S11=39S 95=7X 
 tpg|BK006941.2| 726594 + tpg|BK006941.2| 726503 - INS CCCCTATAGACACCCAGCGGAGCTCCTCCCGAGAAAGGCCCCTTCATCTCTGCCGATTGCTGACGGAAAGCAGTAGCGGAGGTTTGAGTTCTCTACGCCGAGAGTACACTGCCGTAATATCACAATGTTTCGACTAACGGTTACAGTACGTTAAATTAGATACTGCCTATGAA tpg|BK006941.2|:726143-726954 14S79= 87=7X 
 tpg|BK006938.2| 571683 + tpg|BK006938.2| 572011 - INS TTGTTAAGAGTAACTCAAAGTCGGATGAGGAGAAAAGAAAGAAGAACTTTAAAAAGGGTAAACACGGTGGTAAATCTGTAAAAATCGAAAAAACGGAAAATGAAGTTTTAGATGAAAAGAACTCAAAATTATTCAGTGCTTTGTTAACAGGTATCAATCGTGCAT tpg|BK006938.2|:571339-572355 7X23=1X58= 156S1=7X 
 tpg|BK006941.2| 318221 + tpg|BK006941.2| 318397 - INS AATTTATTATCATATATGGTATAAGAAAATGACATGAACATTGAGAAACAACCAATAGATTAATTGGAAGCTGAAATGCAAGGATTAATAACTTGATAAATGGAAGTTAAAAGATAGTATTAATGATGACTAAATATGGATTCTGTTATCCTTGTATAAG tpg|BK006941.2|:317887-318731 7X5=75S 72S8=7X 
 tpg|BK006941.2| 533269 + tpg|BK006941.2| 532848 - INS CCAAAAAGATATAAAAATTTTGTAGAAAAAAAACAACAACGTTGGAAATGGCGAAGACTATCAAAGTTATCAGGAAGAAGGACCCCAAAAAGAAGAACCTATCCGATCCTTTAGCAAAACAAAAACTAGTTTGGAAAATCGGACACGTTTTAAC tpg|BK006941.2|:532526-533591 11S73= 77=7X 
 tpg|BK006938.2| 1429464 + tpg|BK006938.2| 1429621 - INS GTGCACAGACGTAGCCTGAGGAATGGCGTACAAGAAAGGCCATTTGTTCAGTGCTGACATTTTCAGCAGCGCAAATAAGATCACCTTCATTTTCACGACCGGCATCGTCCATAACAATTACAAACTTATTCTGCTTGAAGTGTTCTATAGCTTGATCAATTGGTGTAAACATTTTCGACGTTGCCTTTTCTTCTTTTCCTTTCCTTTTTTTTAGCCTT tpg|BK006938.2|:1429014-1430071 7X6=103S 97S12=7X 
 tpg|BK006941.2| 786540 + tpg|BK006941.2| 786215 - INS GTTCACGTAGGAGAAGGCATTTTACCATACTCCTACAAGGGGCACTAAAGTCCCTGCGCAGTGTATGGGAT tpg|BK006941.2|:786059-786696 7X5=30S 32S4=7X 
 tpg|BK006941.2| 142677 + tpg|BK006941.2| 142437 - INS GGTATTTGCAACGCCGCAGTC tpg|BK006941.2|:142381-142733 7X4=6S 11=7X 
 tpg|BK006938.2| 1134969 + tpg|BK006938.2| 1135080 - INS AAGAGGTGCTTCCTCTTGTCTTTTGCAGCCTCGGCGGTATGGTTTTTTTGCTTCCTTTTTGCCTTTTTATTCTTTTTCCTTCTAGAAGACTTGGATGCTAGTGTAATTCTTTTAGGTTGACCATTACTTTGAGTATCACGCTCCCCAGCAGCAGCAGCTTCTTCATCCTGCTCAGACATTTGTCCTTCATCAGTGCTATTATCTGAATCACGTACGTTATTCATCATAGAGAAGATGTTCTCCCGTTTCTGAATATTACCGGCAGTACTTTTACCACTCGTCATTTTATTCGCATTTGAATTCGATAGCAGCGACT tpg|BK006938.2|:1134323-1135726 7X269= 297=7X 
 tpg|BK006938.2| 417187 + tpg|BK006938.2| 417718 - INS CCGTCTCAAACGTGTATCTGTGGGGGGTAACCATGGCAATAGATGTGGTTGTGGAGCATTCAGCGTGATAGCAAAAGGTGTTAAATTGAATGGCTCCTCAGGACGGTCGTTTGCCTTCCATATTAAAAACTTCGTTCCGTCATCCGTAGGCCCATTCCCTGCTGATGCAGCGGTTCTAGTTTTCTCCAACGAGAGATCGCCATCTTTTACTACTTTCTTGGCAAAAATAGCTTCATTCCAGTGTCCTCCTAG tpg|BK006938.2|:416669-418236 7X230= 126=7X 
 tpg|BK006938.2| 403228 + tpg|BK006938.2| 403236 - INS TAGTGGGGGGTGTATTAGTGCTCGATTTTAAATCCACATAATCATGGAATGAGTTTGTTGACATGTTTGTTTTGAGATCATCCAGTTCTTGCAGAAACAATTTATTATTTTGGTTGTAAAGCTACTTCTATAAACAACTGCAATATTCCTATTCAGACTTCAGTGGGCTGGGTCAAGTAGGCTTCTATAAATTTTGTAGGTTACTATTAATATAGTAGATCTTAAATTCTCTTTAAGCTTGCCTTCACATAAACATCACTATTACTCTTTGCAACCCTTGGTAG tpg|BK006938.2|:402646-403818 7X6=182S 3S264=7X 
 tpg|BK006938.2| 1358326 + tpg|BK006938.2| 1358768 - INS GGTTACCTTAGTGAATTTAATCTATGCTCAAAATCAGTTCTTTTCTTCATAATTAATGAAACTTCATTTTTAGTGAATAGTCCTTTCTCCACCAAGTCATCCATTTCAGGAATACATTGTTCCAAATAGTATCTTGTCTTCGACATTATTAGAAATCGGTGATGTGTGTATCTCTGGTCAATTTCACAATGTTATGCCC tpg|BK006938.2|:1357914-1359180 7X269= 187=7X 
 tpg|BK006938.2| 379504 + tpg|BK006938.2| 379699 - INS CTTTCCGTCTACGATGAACCAAGTGTAAGTCCTTAATACCATTAACAGAATCATCGTTTTTGGTGAAAAGGGACGCGACTTCCACCGCCTTGTCGATATTGTTAGCCCTTAAAAAGTACTTAACCGTTTTACAGTTGATAAATCTATCCTGCAAATCAAGTTGCCTACCTTCCTCCAAAATTCCAGCCGCTGTGTCCATTAGGCCTAAGTGCTTCAGGATACGTGCCTTGAGGATGTAAAACTCAACTAAAGTTGGGGTGTGGTCAAGGGCAGCAT tpg|BK006938.2|:378938-380265 7X191= 242=7X 
 tpg|BK006938.2| 633052 + tpg|BK006938.2| 633138 - INS TCCTATGTTTCAAGATTATTATAAACAGAAACCTCGATCGAGAGATTATTTTGAATTTGGTACCATTGGAGGTTCTGCCTCAACTAACGGTTTTGTTTCTTTTTGGGTGGCGGTTATTCTTTATCAGTCATTGGTTCCGATCTCTTTATATATTTCTGTGGAAATTATTAAGACAGCACAGGCTATTTTCATTTACACTGATGTTTTGTTGTATAATGCCAAGCTAGACTATCCATGTACACCAAAGTCGTGGAACATCTCCGATGATTTGGGTCAAATTGAGTATATTTTTTCAGATAAAACAGGCACCTTGACACAAAATGTGATGGAATTCAAAAAATGTACTATTAACGGTGTGTCTTATGG tpg|BK006938.2|:632306-633884 7X203= 344=7X 
 tpg|BK006938.2| 707391 + tpg|BK006938.2| 707526 - INS TGTGGAGGGATGTGGAAGAAATTCGTGAAGTTTGGAACAGAAGGGAGGGGTGGTATAAAGAATGCTCAAATTTCTCTTTCTTTGCTCCTCATTGCTCCGCAGAAGCTGAGTTCCAAGCTCTAAGAAGATCGTTTAGTAAGTACATTGCAACCATTACAGGTGTCAGAGAAATAGAAATTCCAAGCGGAAGATCTGCCTTTGTGTGTTTAACCTTTGATGACTTAACTGAACAAACTGAGAATTTGACTCCAATCTGTTATGGTTGTGAGGCTGTAGAGGTCAGAGTAGACCATTTGGCTAATTACTCTGCTGATTTCGTGAGTAAACAGTTATCTATATTGCGTAAAGCCACTGACAGTATTCCTATCATTTTTACTG tpg|BK006938.2|:706621-708296 7X341= 367=7X 
 tpg|BK006938.2| 1035799 + tpg|BK006938.2| 1036421 - INS AAAATAGGACCTTTCTTAAATGATCAGGAGATAAAGGTTTCAAAAAGGCCATTGATTTTGCAAAAATCCTTAATTGCTTTAGAAGGAGGTTCGGAAAGAACTGAAGGTTCCCAAGGAAACTTTGATAAGAAAATGAATACTTATAAAAACTTACTAAGTGAGTCCGGCGCCTTTGTTCACGGGTTCAGAAGTGCAGGAAGTGCTGCCATGAACATATGCTACGTAGCGAGCGGCATGCTTGATGCTTATTGGG tpg|BK006938.2|:1035279-1036941 7X7=223S 238=7X 
 tpg|BK006938.2| 594400 + tpg|BK006938.2| 594983 - INS TCCCTGGAAGTCTCAGCTGATTCATTTAAATACTATCAATTTCCGTGTACTTTCGGAGATCTTTCAGTCAGCTTTTCCTTCATCTTTTTCAGTCTAATCTAAGGAAGAAGAAAAGCACTTCAATACGAATAGCTACCAACGTACCCAGTTCACGTTGAACAAGCAATAGAAAACCAAAATA tpg|BK006938.2|:594024-595359 7X5=85S 86S5=7X 
 tpg|BK006938.2| 1037326 + tpg|BK006938.2| 1037747 - INS TGTATAACGTATATTGGTGATCGTCATTTTATGCATTGTTTTCTTCTCTAAGAATAACATATTACATCAGGAATTGATCAAATTTCTAGAGACATTTGGCATTCCAAGCGATGGTTCAAAGATTGCTATACTGAACATTACTATTGAAGATTTGATAAAAAGTTTAGAAAAGCGCGAATATATAGTCAGATTGGAGGAGAAATCCGATACCGACGGGGAAGTGATATCATACAGGATAGGTAGAAGAACTCAGGCTGAGCTTGGACTAGAGTCTCTTGAAAAATTGGTGCAAGAAATCATGGGCCTTGAAAAGGAGCAGACTAAAAGTTTGCACGATGATATAATAAAAAGCATTGGCGATTCATATTCTATATAGCATTGCATAGGTGTCCAT tpg|BK006938.2|:1036524-1038549 7X4=156S 370=7X 
 tpg|BK006938.2| 396228 + tpg|BK006938.2| 396153 - INS ATTAGATTTGAAGATGCGGACCAATTATTAGAAGCACAGGAAAACGAAAACAAAAAGAAAAAGAAACCGAAGTCTTTTAAGGATCCAACTTTCTTTTTAAGTCACTATGCGCCAGCTGGTGACATACAAGATAAACAATTACAGATAACCAATGGGTTCGCTAATGATGCTGCTCAAGCGGCTTACGATTTAAATAGCGATGATAA tpg|BK006938.2|:395727-396654 12S162=19S 15S5=7X 
 tpg|BK006938.2| 839868 + tpg|BK006938.2| 840580 - INS GCGTGTGCTTTAGGCTTTCTTCACTGTTACAAATAATTTGCGGAAGTTTCTAAAATCTTTGTTGACCTTTTGGCATCCAAAAACAGCAATTTGGCTTCATTAACGTCATTAACAACAATTTCCTTACGATTGCTTGTTTGTGCTAGGATACCACATGGTGCCAATAATTGTAAAGCGTAACGTAACGAAGTTTCTGTACCCATCGTGGCTAAAAGGTCCAATGCGCTACTTTCTACTTGCAATCTTTCAACGGTAGCTCTTCTCTCTATAATGGTACGGATCTCGTCCTTGTCATATGGTAATGTACGAACAATTAACAATCTATCGATCAAATCAGGTGGCACACCATGTGGTGATATCACATCCTCAGTGCCACGGACTGTAGTCATGCCCCTATTAGAAGC tpg|BK006938.2|:839046-841402 7X50=1X209= 202=7X 
 tpg|BK006938.2| 1492129 + tpg|BK006938.2| 1492128 - INS GTATAACTCTTTAGATCCCAAACTGATTGCCAAGCTATTGAAAAACATAAATAAAAGAGCGAAGGACGAAAACAACACTCCATTATTTGCAGAAATAGAAGGCGCTTCTGGTACCTGGGTAGGTGGCAACAAGCAAGGCATATACGATCTACCACCGTTAGACGATGAAGATGTAGACGTTGCCTTAGAAATTAGGCCTATGTTAGGCAAAGATGCAAAACATGTT tpg|BK006938.2|:1491662-1492595 7X4=109S 107S6=7X 
 tpg|BK006938.2| 750096 + tpg|BK006938.2| 749730 - INS CTCTTGTTGTTAGCAGAGTTGGACGTAGCTGAACTAACTCTACTCTTTGGAGTGAAGGGCGTAATAAATTTGGTTTTTGAACTGAGGTTTTCATTTGGATTCGAGCGAATTTTCTTTGGTGAAATGAGGGAGTCATTGAAACCTTCGTTCAATTCCTGGAAACATAGTGGTCCTACAG tpg|BK006938.2|:749360-750466 7X276= 89=7X 
 tpg|BK006938.2| 1504187 + tpg|BK006938.2| 1504664 - INS TGTTGGTAATACTTTCGCCTAAAGCGGCAACGGTGATAGCAGATAATACAAAAGCGGAAGACAATTTCATTTTCGGGTATTGTATTGTTATTACTATTATTATTCAGGCGAACAAAAGGACTTTCTGAAAATAAACACGGCATTAGGAATATAGAAAAGTTAGATAATCATTAGTTTAAATAGTGCAAAAACTTCACTTCAAAAATGGTATACGAGTGTCATATTATATTAGATATTCATTTTTTTGCACCCTTTCCTAGAACTCGCGTATTGAGCCCTGAGGTGTCTGTCATTACATTATGCCAAATGTGCGACAGCGCGGTTTGGAACAAACAGGGTGCGGAACAGGGT tpg|BK006938.2|:1503471-1505380 7X158= 176=7X 
 tpg|BK006938.2| 843102 + tpg|BK006938.2| 843504 - INS GGCATTGTTTGCCCAAATGAAGGGTTCGATTGCGAGACTTTGTTGGCATCGTTTTGTGGTGTAATTCCGAATGAAAACCCTTTATTACCAAAAGAAGATTGAAAGTTGCCATTGGTATTTTTATTGAGGTTAGAAGCAGAACCAAAGGTGCCCCCAGAACCTCCGCTAAAAGGAGATTGATTATTCGTCGTTCCGAATGCGCTACTGCCCACGTTATTGTTGTTGTTAGCTTTGGAGGTTGTAGTACCAAACGGCGAAGAACCAGCGCCTGCTC tpg|BK006938.2|:842540-844066 7X236=15S 2S1=228S 
 tpg|BK006938.2| 897223 + tpg|BK006938.2| 897211 - INS CCTTTAATGGCTTATGATTTTTGTCAGTTCTTGAAATGTTTCGTCCATATTAAATTCGATTTGTCTATAAAGGAAAAAGATGTTGAAACCATTTATATTCCCGACAATGAGTCAAAATGGGCCAGTGAATCGATAATATGTAATGGGCATGTTGTGCAAAAGCAAAATTTTTATGATTTTAGAAACTTTTATTACAGTTTCACGTATGGACACTTACACTC tpg|BK006938.2|:896755-897679 7X2=1I39=1X76=46S 1S1=148S 
 tpg|BK006938.2| 159200 + tpg|BK006938.2| 159753 - INS CATCAAAGTTGTCCTCGTGTGCATCATATACCACCTTATATGATTGTTGGTATTGTGTGGCGAATAAGTCCTGGTTCCAGGCAAAACCTTGACTTTGAGATACAGATATTTTAAAATTTGGCCTTATTTCTGCACTATATGTAAATACCGAA tpg|BK006938.2|:158882-160071 7X5=71S 70S6=7X 
 tpg|BK006938.2| 589834 + tpg|BK006938.2| 589214 - INS CCAGATACCATCTCTCTGATGAAAAGACCTGAACATAGCTCTGGACAATTGATCAAACGAAAGCTGATAATTTCTTCTGAAGCTCTTTCGTTTGGTGGGAAACCTTGGCTTTCCAAGTTCAAAATCTGCTTTAAATCTTCAATGATTAAGGGTCTAATATACATATGAAGCGGTAGCGTGCTACTTGAGG tpg|BK006938.2|:588820-590228 7X4=182S 179=7X 
 tpg|BK006938.2| 596193 + tpg|BK006938.2| 596536 - INS GGGTGATGACTTATGTTATGAAAAGATCGGCTTCTTACACCGGCGCAAAGGTTTGAAACACCCTTTTTAACGAAATGGTTATGACTAGACAGACATCTTACGTCTTACTCCTTCATGCTTTATTTTTTTCTTTGTATTGTATTTGAACAGTCAATATGTGGTGTTGCGACGAAGGCATATATATAATAGTCTCAACCCACCATTTTCGAAGATTTACATACACATTATATTTTTATAAACTTCCAATATGTAATAACTTTATATGATATGTAACTTCTCACTATTATCCTTACTATTAAACGGTTTTTAATAAATATCATTGTTCTTTGTTTTATTAATGAGAAAAAGAAATTTAATACAATGTCCGGCGGGAAGAAAAAAAATCGATGAATTAATTGAAAAAAAGTATCTTTATCATGTGAACTGAGGAGAAGAACGGCATCTCGAAAAGAGCACGTCGAAACAGCGGTAGGT tpg|BK006938.2|:595231-597498 7X268= 460=7X 
 tpg|BK006938.2| 1050774 + tpg|BK006938.2| 1051193 - INS GCCTGGACCCTAGACAACTGTCGACGTGTAAAGGAAGTTTATATTTTTGTGCTATTTTACCCAATCCTTCAATATCATCGGCAATACCATGAGGAAAGTTTGGAGCGGAACCGACCAGTAAAATTGTGTTCTTATTGATGAATTTTTTCACTTTTCCCAGGTCCACTTGATATGTCGTTGGATCTAGCTCCACGTGGCGTAGCTTCATGCCAAAGTAATAAGCAGCTTTGTCAAACCCAGCATGTGCAGTTACGGGAGCAATTATTTCTGGTTCGGTGATTCCACGATGATGAAGGGCATACATTTTAGCGCTCAGACATGCTAAAAGC tpg|BK006938.2|:1050102-1051865 7X399= 309=7X 
 tpg|BK006938.2| 1043006 + tpg|BK006938.2| 1043037 - INS ATATTACATCAACATTCTGTCACCTTGTTGATGCACAGAAAAAAAGACACTTTATTATTGTTGAATAACATTGTCTGTGGTATATATATATATACTATGATATTACAGTTTTTAAGACATTAATGTATTAACAGCCCATTTTACGCTTAATGTCCTCAAATCGGTATAGGTTTGTCC tpg|BK006938.2|:1042638-1043405 7X157= 89=7X 
 tpg|BK006938.2| 511144 + tpg|BK006938.2| 511075 - INS TATCTCTTAACGAGGCTAGTACATTATTCTTGCTCTCTAGGGATTCTATTTCATCCAAAGGTACATTCTTGCCGTTATCTGTAATCGGTTTAGGGTCCGTGGTGTCTTCACTTAAATTTTGTCGTACTTTTTTCTTCTTCTCAGCCTTGCATGACGAATGCTGACGCTTGCGAGCATTAGTATGATCATTATCGAGGCTAGTACTGTGCTTCCTAAATTCTTTTACTCTTTGAGCATTTGAGGTTCTTCTTTTCTTATTTTTTGGGTTTAAAACGTAAACGCACTGACGATTCAATCTTGCGCACTGCCAACAAGTCGGTTTAGTTT tpg|BK006938.2|:510407-511812 7X120=1X167= 13S146=1X147=7X 
 tpg|BK006938.2| 1138704 + tpg|BK006938.2| 1138928 - INS TATTGTAAGCCCCAGACTGACGTGTGTAACTCTGCTTAAATTGTTCAAAAAAAACAATCAAGTTAACCGGGTTGACTTGGATTTCTTGAACTTGGTGTTTACGCTTAATGACAAAGATTTAACTTCTTATCATGCCGAGGAAATCTCAAAACTGACGTGTGTAAAAAACTTCGTTGAAGAAGTCAATAAATTGAGGGAAACCAATAAACAGCTTCAGGAGGAGTTTGGAGAGGCGTCTTTTTTAAATTTTCAAGATGCAAATCAATATTTCAAGTATTCTAATAAGCAGAAACTTGAAGGGACAGTTGACATGCTAAACTTTCTAAAGATGGTAAATAAAC tpg|BK006938.2|:1138008-1139624 7X310= 7S313=7X 
 tpg|BK006938.2| 501213 + tpg|BK006938.2| 501385 - INS GTGTGGTTCTCCTGTTCTCCTGTTCTCAGGGCTGATTCCTTCCTTCAATATCCACTGTGAGTTTAAATGCAAACAAAAATAGAGTGAATAAAAAAAGCTTTCGGCCCGGAATTGGTTAACCCGACTTACCAATATTATGTCAGAAAAGAGGCTACAGCTGAAACTAAGGTGAGGTGGTAAGAAATGCTCTCTATTGAAAAGTATGCATGAAGTGGAGG tpg|BK006938.2|:500763-501835 7X4=388S 10S195=7X 
 tpg|BK006938.2| 356469 + tpg|BK006938.2| 356754 - INS CAAGAGCGTTGGCTTTACTACCGGTTTCCTTTTCATTTTTCAATTATATATGTTTTATTTGTTGAAGTTGTAGCTTGTCTTGTGCTGATAATATTTTGTTTGTATAGTCAACAAAATATTTGGACAGAAGAAAAGAGTTAGCGAATGTAAAGTAGTTTGCACACTTGATGAACGTTATCAAAGTCAAAGAGGTGAGAAC tpg|BK006938.2|:356057-357166 7X162= 12S169=7X 
 tpg|BK006938.2| 614873 + tpg|BK006938.2| 614875 - INS ATTTACCATGTCATTCATAACCGTCATCATCATCAGTTTGACTTTCTGGCAAGCTGGTCAGGGTATTAACAGCAGATATCGGAGAGGTTGATGAAACCGAACTTTTTATTGTTGAAGGAACTGAAGTGTTCAGCTCCAAGCTATTTACACCGTAGCCTGTATCATTGGGAGGAATATGTA tpg|BK006938.2|:614499-615249 7X12=78S 86S4=7X 
 tpg|BK006938.2| 1095489 + tpg|BK006938.2| 1095127 - INS GTTCTCCTTGTGAATTAGGTACACAGAATATTCATGAAGTTTTTTTTGAGGATAAAAGAATCCCCAAAAAATGAGATTGGTAAATCTTGTTGGAATAAAAATCCACTATCGTCTATCAACTAATAGTTATATTATCAATATATTATCATATACGGTGTTAAGATGATGACATAAGTTATGAGAAGCTGTCATCGATGTTAGAG tpg|BK006938.2|:1094707-1095909 7X197= 191=7X 
 tpg|BK006946.2| 773655 + tpg|BK006946.2| 774127 - INS TCTCACAGTGGGGTATACGAGCACGCTTGTAAGGGGGATGGGGGCTAAGAAGTCATTCACTTTCTTTTCCCTTCGCGGTCCGGACCCGGGACCCCTCCTCTCCCCGCACGATTTCTTCCTTTCATATCTTCCTTTTATTCCTATCCCGTTGAAGCAACCGCACTATGACTAAATGGTGCTGGACATCTCCATGGCTGTGACTTGTGTGTATCTCACAGTGGTAACGGCACCGTGGCTCGGAAACGGTTCCTTCGTGACAATTCTAGAACAGGGGCTACAG tpg|BK006946.2|:773081-774701 7X4=202S 1S262=7X 
 tpg|BK006938.2| 971059 + tpg|BK006938.2| 971520 - INS GCCTTGATTATCACCACAAGGACAAGTGGCAACTACTGTGTGTATACAGATTAAGCTTTTACAAAGGTAATGAAATTTTTTCATACTCGAGAGAAAAATATGTGACACATGTGTGTATTACCCGCAGTAACTCTCGAAGATTACATTTGAATAATATCAATACTTCCAGACCAATAGCTTTATTGTATTGCCAGGGCACTTGGTACATGTAACATTCATCCAGTTTATTTGATACCAAAAATCTTTTATTTTAATTCTTCTATTTACAAAAGAGAAATGTGTATGTTTATATATGTATTTTCTTGGGAATTTATTATTCATAAACCGCTTGTGCAGTTACTTTTCAGCTTCCTCTTCAACAACTTCGCCTTCTTCATGATTTGGTAGCACGACAAGCTTAGTATCTTTAACCACCACTCTAACAGTTTCGCCGTTTCTAATTTGACCTTTTAATAAGAAAGTTGCCATGGAGTTCAAAATCTGTCTATGAATTAATCTATTCAATGGCCTTGCAC tpg|BK006938.2|:970015-972564 7X158= 17S466=7X 
 tpg|BK006938.2| 1221220 + tpg|BK006938.2| 1221967 - INS TTGCCCCATATCAAAAGTTGTAATGAAAATATAGCCAACAATGAAACTGCTAATTTAGCTCTATTTGTTAGCGTGGAAATTTGAAATTTATTTTTAATCTATAAATGCAGCAGCCCAAACCGAAACAAAAGAATAAGTGAGTTGAACAGAGTAAGCAACGGGCCGATATAGAACTGAAAAAGTCAACGTACCCAGAAAGCAATTAACTGCGACACAAATAGATGTCAATGTCCAAAAAGGATAGATAAACAAGATTACGATCCAAGGC tpg|BK006938.2|:1220670-1222517 7X166= 252=7X 
 tpg|BK006938.2| 435941 + tpg|BK006938.2| 436655 - INS TATTCTTTTTTCTTTTGCGGTGGTAATTACGGGAATTTAGTGATGTTGGAACGAGAGTAATTAATAGTGACATGAGTTGCTATGGTAACAATCTAATGCTTACACCGTATATTAATGTACACCTCGTATACGTTTAAGTGTGATTGCACCTATTGCAGAAGGAATGTTAAACGAGAAGCTCAGACAATACTGAAGCTGTGCTAAAGATCTATTAATTGAACATGATATGGTAGGTACATATATGAGGAATATGAGTCGTCACATCAATGT tpg|BK006938.2|:435387-437209 7X104=31S 1=168S 
 tpg|BK006938.2| 1324245 + tpg|BK006938.2| 1324614 - INS TATAAGGTGGAACATACTGCCCTGGGATGGAACCAGCTCCGCCAACTTGGCCTGCCTTCTCTTCACTGGCGGCCTCGACACCGCCTTCATTAGTGGCTGGGTCTTCTAATGCTGAAAGTTCACTTAAAATTGTCTTGAATGGACAGTTCATGGTCATATGGTCGTTACCACATAATCTAC tpg|BK006938.2|:1323871-1324988 7X153= 90=7X 
 tpg|BK006946.2| 910958 + tpg|BK006946.2| 911095 - INS GTACCTTATAATTGATCGGCGCCCATCTTCATTGCATCTTCTCTTTTTCTCGAAGAACGAGAAATAACATACGTCTCTGCCCCCATGGCTTTGGAAATCAATGTACCCATACTGCCGATACCACCAAGACCAACTATACCAACTTTTTTACCTGGACCGCAACCGTTACGAACCAATGGAGAGTACACAGTCAAACCACCACATAATAGTGGAGCAGCCAAATGTGATGGAATATTCTCTGGGATAGGCACCACAAAATGTTCATGAACTCTGACGTAGTTTGCATAGCCACCCTGCGACACATAGCCGTCTTCATAAGGCTGACTGTATGTGGTAACAAACTTGGTGCAGTATGGTTCATTATCATTCTTACAA tpg|BK006946.2|:910194-911859 7X273= 352=7X 
 tpg|BK006938.2| 43276 + tpg|BK006938.2| 43879 - INS ATCGAGGAGTTATCAAGAAAAGCGTTTGTTAGTAGTAGTTTGCGACAGTGGAGATGGCAGCTGCACCATGGTATATTAGACAGCGTGACACGGATTTATTGGGTAAATTCAAGTTCATACAGAATCAAGAAGACGGCAGATTAAGGGAAGCTACAAACGGAACGGTGAATTCACGATGGT tpg|BK006938.2|:42902-44253 7X5=85S 84S6=7X 
 tpg|BK006946.2| 67397 + tpg|BK006946.2| 68060 - INS CCATAAATGTAATCCGATTCAACTCGAAGGGTGACGTACTGGCGTCTGCGGGCGATGACGGCCAAGTGCTGCTATGGAAGCAAGAAGATCCAAATACACAGCAAGAATCTGTGGTCAGACCATTCGGAATGGATGCGGAGACTAGTGAAGCAGACGAGAACAAGGAGAAATGGGTTGTGTGGAAACGGCTGCGTGGTGGTAGCGGTGCTACTGCGGCGGCAGAGATTTACGATCTAGCGTGGTCACCTGATAACAGGAACATAGTGGTGGCATGTATGGACAATTCGATACGACTGTTCGATGTTGGAG tpg|BK006946.2|:66765-68692 7X182=49S 7S1=185S 
 tpg|BK006938.2| 870730 + tpg|BK006938.2| 870652 - INS GCAACAGGGTGTGTGGGGCTTCCGCAGTGTGTGGCTAAGCGGCTTTAAGAGGATACGAAATGTCAAAAAACGAGAAAATTCGATTATATCTGTACGAACTTTTCTTTGCGCTTACTGCCTGTTTACTTTGCTTTGCCTTCTACTGTTTTTTTTTGCTCGAGGCCGATGGTGAACTGCAACGTTATATAAACTAAAGTGCCAGAATAAAAATAAAGAAAGGCAAAGGGAGACTATCCGTCTTCGAAACAAGTCAAAAGAGCGAAAACTAATGAGCCAACAACAAGGTTACTACCAACAAGGACCCCCACAGCAAGGTTATTATCAACAAGGTCCACCACAACAAGGTTATTATCAACAAGGTCCACCGCAACAGGGTTATCCTCAGC tpg|BK006938.2|:869866-871516 7X283= 362=7X 
 tpg|BK006938.2| 111549 + tpg|BK006938.2| 110909 - INS GGATGGCTGAAGCGGCAAATCTTGCCGCATCGCACATTCTAAAGAACAAAAGGAGGAGGAACTGTCAATTATTCTATAATCTGGGGAAATTCAGTCATACTGAGAAAAACTAGACAATAGTCCTATCCTCGGCAAATTGCATTGATAGTACTTACACATCGAGAGATCATAGGACAGATAAGAAG tpg|BK006938.2|:110525-111933 7X4=222S 9S165=7X 
 tpg|BK006946.2| 500739 + tpg|BK006946.2| 500158 - INS TAGTAAATCCGTACATTTTGTCGTTACCGGCAGAAATGATGGTGACAGAGTCATCATCAGCTTTTTCGTTTGGAACAACTCTGACTTGGGAAACCCAGTCATTGTGACCCAACAAAGTGGCCAAACATTGACCTGTGATGGTCCAGACCTTGATGGTCTTGTCACGGGAACCAGAGATAATCATGGAAGCCTTCTTGTCAATGTCAACGGACATAACATCGGACTTGTGACCGACGAATCTTTGGTAGGTTTCACCGGTGGCAACATCCCATAATCTCAAGGTCTTGTCCCAAGAAGCAGACAAAGCGTAAGCACCGTCAGCAGTCAAAGTACAGTCTTGGACAATGTGACTGTGACCCTTGAAAGATCTAACTGGGACACCAAACTTTTGGTCGTCACCAGTCAACTTCCAGGAGATCAAAGTCTTATCACGGGAAGCGGACAACAATAGGTTTGGTTGACCAGCAGAAG tpg|BK006946.2|:499202-501695 7X4=1X5=299S 120=1X336=7X 
 tpg|BK006938.2| 1076186 + tpg|BK006938.2| 1076933 - INS CTACGACAATGAAATCAACAATGATAAAAAGGATAACGCAGATGATAAATACATTAAACCGCTTCAATCAGAGATACGCTTTTACAATAACGGCCAGAGATGTGGGCTATTGGGCCATGATCTTCGGTTACCTGAATGGGGCCGCTTTGAGCAAGAAGTCCTATGTATGGAGTACCCAGTAATACCAAGAACCACTTTTCTAATAGACTCAGTACAACTACCAGTCGATTTCCAAGTCCCAATGATAGAATATTATATCGGCAAAATAAGTTCTTCAGCAGAATTCAATCATACCT tpg|BK006938.2|:1075580-1077539 7X385= 278=7X 
 tpg|BK006938.2| 1500795 + tpg|BK006938.2| 1500846 - INS CACAAACTTGTTCGTGGAGACCAAATGTATTCTTCACTATTAACCTCTAGCTAAAGCAGATAAAAGATAAAGATTATAAACTTTGGTTATTGGAAGACCCATCTCAGACATGTGTTTCCCCAATATCCAAATATTTCAACGTATTAACAATGAGGTACATCCCTCGTACTCAATAACGCCTCCTAAAGTTCCTTACATCTATATAGT tpg|BK006938.2|:1500367-1501274 21S15=1X39=34S 98S6=7X 
 tpg|BK006938.2| 1309828 + tpg|BK006938.2| 1310243 - INS AAGGCATACATCATCATTATCAGTTGTCAAGAAAAAAAAAAACCAGCAGAAAAAAAATGCCACGAAGTCAACCGAGGACTTACATCCTCCACAAGTCGACACATCCTCAATAGCGGTGAAAAAGATTGTTCCCATGGTAGACTCTTCTAAGG tpg|BK006938.2|:1309510-1310561 7X5=208S 133=7X 
 tpg|BK006938.2| 1006721 + tpg|BK006938.2| 1007289 - INS CTTTGTTAGAGGTATATTGACTTTCTTTATTTGGTGTTTTATTTTAAACATCTCGGCTAATCCTCCCGTCGCTTTCACCGCAAATACTAAGGCTGATAATTTTTTTATTTGCTTACAAACTGCTACTTCTGTTGTCATCGTCGCATGCCCATGTGCATTGGGACTTGCCACGCCGACTGCTATAATGGTGGGTACAGGGGTTGGAGCTCAGAATGGTGTCTTAATAAAGGGCGGAGAAGTATTGGAAAAATTCAATAGTATTACTACTTTTGTTTTTGATAAAACAGGTACCTTAACTACAGGTTTTATGGTTGTGAAAAAGTTCCTTAAAGATTCAAATTGGGTTGGAAACGTGGATGAAGACGAAGTTCTCGCCTGTATAAAAGCAACGGAATCCATTAGTGACCATCCAGTTTCGAAAGCAATTATACGTTATTGTGATGGTTTGAACTGTAATAAGG tpg|BK006938.2|:1005785-1008225 7X200= 447=7X 
 tpg|BK006938.2| 162101 + tpg|BK006938.2| 162241 - INS AGATAGTATTACAATTGTTGTTGGAGATTGCTTTCTTTTGTCCCAAAATCTCCGGATGGTTGACACACCATCTATCGAATTCCTTCCATAAGTCAAATACTTTCGGATGTTGTAAATAAGAAGTAAGAATAAACCCATCATCTCTCGCTTGACGTGGTAAGGTAACACGGATATGCCATGTTGAATACAGGGAAACAAGAACAAAGTCGTCGTTACCAATAACGTCATGAATATCCTTGTCCAATTGCACCATTGCAC tpg|BK006938.2|:161571-162771 10S47=79S 125S4=7X 
 tpg|BK006938.2| 523483 + tpg|BK006938.2| 523482 - INS CCTGTTCTGTGATCTCTGGAATTCTCTTGCACCAATCTCAAGGCGATTTGAAGAGAGGATGGTGACTTGGTTAACAATTTCGTTTTGATTTCTTGTGCGAAAGCCTTACCTTCCGCAGAACCTTCATATTGACGTAAGTTATTCATTATGTCTTCAATAGTACCATTTTTAGACAAGTTAAAACAGGCTTCAAT tpg|BK006938.2|:523080-523885 132S147= 97=7X 
 tpg|BK006938.2| 23964 + tpg|BK006938.2| 23198 - INS GTTACAGATATGTGCTACTCCTTGTGGGGTTAAAAAATGCTTCATGTACGGAAACCAATTGTATTGCAAGTACCACTTTCTCAAGTATTTTTCGAAACGTTGCAAAGGGTGCGAGTTCCCAATATCGGATCAATATATCGAGTTTCCTAAAGGTGAAGAAATACATTGT tpg|BK006938.2|:22846-24316 7X7=306S 85=7X 
 tpg|BK006946.2| 777292 + tpg|BK006946.2| 777254 - INS TTACCTTCGGTCTCTACGTCAAGTAAATATATGTCAATATATCGATGTGTCGGCAGACTTGCTGGCTTGCGCGAGTTAATGAAGTAATAGAACAAGCTTTCTGTAATCATCCCGTCACTTATGCTTTTGTACATATCGTGTCATACTGCGACTGTCTCAAGGAAATACCATGATAAAATATCTCTTACAATCGAAAAATCTAGCACGTGGGAGGGTAAGCATAAACTACCCAGAAACGCATGTATGGACTGCATTTGCTTCCTGACCAAAATAAGTATTATCGTCATATAAAAAACGTGCATAGTATATGTAACATCAATGATGCTGGGCGTTGTTTGCCATTTTGTATTTACTATGGCAGTGTATTTTGTAACGAGCACGTGATTTACAGGGCGCAGAAATGTTGAAAATTTAGAAAAAAGTAAGATAAGCAATATCAGTGGCACCATTGAGCTAGTCTCTAACAGCGGGGTGAGAAGC tpg|BK006946.2|:776280-778266 7X295= 465=7X 
 tpg|BK006938.2| 1523306 + tpg|BK006938.2| 1522702 - INS AAAGGTATATGTTTCACGTAAAAGGGTTCTTCGAAGGCACATGGCGCCCCTATAACGTCGATCTTACATTGCACGCATACGAATACACATTGGCGCCGCAAAACATATCTTCATATACGAAGTTTGTGACGAATTCACGAATCGTTCAAGGACAGGTGCATTTCTATAGTTACGGTGGATAAGGT tpg|BK006938.2|:1522318-1523690 7X220= 3S171=7X 
 tpg|BK006938.2| 728041 + tpg|BK006938.2| 727367 - INS ATCGTGTAAATCCAAAGTTTTTTTTCTTGCAAAGGTTAACTAAATCTCTGATACCGAAGGTTATCATGAAAATTGCTGATAGATTTAGGATCACACCGTCGATGAAGCATTGAGTAAAGTCACCGTAAAAGGATATAGGTCCAAACCCTTCAGGAGATCTACAGAGCTTGCAGGCCCATGAAACAAGATTACCAGCCATTTTCTTGTTCTTTACGGTAGTACGATACCCCTAATTTATTCTCAAACTGTTAATTGAAAAATTGTAGGTTGTAAACCAGCTTCCACATAGCAGATGATCACAAGAGGTTATCGCACCTTTTATAGC tpg|BK006938.2|:726703-728705 7X5=304S 9S306=7X 
 tpg|BK006946.2| 771399 + tpg|BK006946.2| 771567 - INS GGAATGCCGATTGGTTCAATTCCAAAATTCTCTATTTGTTGCAAGAGCGTTTTCTTTCGAATTATTGAATTCGTCAAAATTGCCCGGATGCTTTGAAATTGTTAGCAGTATCCATGAAAGCATTGAGAACGATTCCGCCCCTAAGTCAGTTAAAGACTATTGGGAACACCCCCAGGCTTACAAACCAGGTGTACCGCTGGTAGCCTTCAAATTGTCCAAGAAATTCCACGAAGAATATCCAGAAG tpg|BK006946.2|:770895-772071 23S106= 16=114S 
 tpg|BK006938.2| 438559 + tpg|BK006938.2| 438411 - INS GGTTAAGGCGAAAGATTAGAAATCTTTTGGGCTTTGCCCGCGCAGGTTCGAGTCCTGCAGTTGTCGTCATTTTTATATTCCCAATATTTTTATCACTCCGGGTAACGAGTTATTAACGGTTTTTCTCCGGTGGCAAATGTCTCTTTTCTTTTACCTAAAAGAAGGTTAATGTGAATATTAGTGAAT tpg|BK006938.2|:438025-438945 7X4=89S 89S4=7X 
 tpg|BK006938.2| 168295 + tpg|BK006938.2| 168347 - INS ATCATCAAGTGTCCAAGGACTCGTTAATTGAGCTGGCTGAAAAATCATATGATAGCGCAGATTTCTTCGAAATCATGGATATGCTGGACAAAAGACTTAACGACAAGGGCAAATACTGGAGGCATATCGCAAAGGCATTGACAGTAATAGAT tpg|BK006938.2|:167977-168665 7X9=67S 70S6=7X 
 tpg|BK006938.2| 264429 + tpg|BK006938.2| 264376 - INS CTCTCTCATTGTAATTGTTTAGCACAATTTCGTTCTCCCTGACAGAGTCCTTGTACAGCGCCAGGTCTCCCGAATCAATGTTCTCCAAGTCGTCGCTGTCGTCAGCTTCAAGACGGTCGTCAGCACCCTCCAACTTAGCTATGTATTTACCCAAGCGGGCGTTAGACCTCTGCAAATG tpg|BK006938.2|:264006-264799 7X133=22S 1S1=204S 
 tpg|BK006938.2| 603439 + tpg|BK006938.2| 604172 - INS CAGGGGCTATATGACGAAGATGAGCCCCCCTTATTGAAGTACACACGAATTAGTCAACTCCCGAAGAACTTTTTTCAACGAGACTCGATCTCTTCATGTTTATTTGGTGATACTTTTTTTGCATTTGGTACACACTCAGGCATTCTACACTTAACTACATGCGCGTTCGAACCCATTAAAACCATCAAATGCCATAGATCTTCGATACTTTGTATTAACACTGACGGAAAATATTTTGCTACGGGATCTATTGACGGGACAGTGATTATCGGATCGATGGATGATCCACAAAACATTACACAATACGATTTCAAAAGACCTATAAACTCTGTAGCGT tpg|BK006938.2|:602751-604860 7X621= 327=7X 
 tpg|BK006946.2| 237004 + tpg|BK006946.2| 237070 - INS GTCTTGCCTTTTGGTCATGGACCACCGAGATTTTCCAACTTTGACATTGAAGATCTTTTTCAAGCAAAGTTTACCAAGTTTATTAAGTTCAAACTGTTTTGGGAGATAAATAAAAATCCAAGTATTTCTACTTTGAAATCGGGGTCAATCTTTGATCAAAATTTCAAACGTGACTCGAAGGTAGCATTTGTCGAGTTATATACATCCCGTGATATGGACAAAATTTTGAACTATTGGACCACTCCTTTGAAGGAAATTTACCACATTACAACAGCGCCCGCAGAATTCGAAGATTTTAAGGATTACAGCAC tpg|BK006946.2|:236368-237706 7X188=1I195= 1S291=7X 
 tpg|BK006938.2| 1126645 + tpg|BK006938.2| 1127019 - INS CATTGATTCATTTACAGGCAGCTTTACTTTTTAACGGCGAACTTTCTCTGCTTTCACTAGACTTTGCTCTAGTCAACTGGTTCTTTTGGTCCTTTAATTGGGTAACGATGCTGTCCAAATTCAAATCGTTTTCATTCAAAACCATTCTCCATACAGGAAGTAGCTCGTATATTGTGTACAACGAGTCTTCCTGTG tpg|BK006938.2|:1126241-1127423 7X179= 6S177=7X 
 tpg|BK006938.2| 295817 + tpg|BK006938.2| 295991 - INS AATAATAAGAATAGGTGGATTAAGTTACAAGTGTTTTTGTCCTCCTACTTAATCAGAACAGAGCACGGGAATAGTGATCTCTTTCAATAGCGAAAGGAGGGAAAAATAGCCCTGCAATATATAAAGGAAGAAGTTAACACCGTATTAAAAGG tpg|BK006938.2|:295499-296309 7X5=71S 71S5=7X 
 tpg|BK006938.2| 154965 + tpg|BK006938.2| 155134 - INS AAGAAGACGGGGACGTTTCTCCAACCTAATACGGATAAGTTGAAGGATGCAGCTAAATCCTCGAAAATCTTCTGACACTTAATTAAATTTTTCTTGTTATTTTTTTCGTTCTTCTTGAAGAAGACGTTACCTACGGCGTATTTGCCCATCTCAGGTATGTCTAGATCAAGATCTAACTTGAATTCTCTTTTCATAAATTCGTGAGGAATACCTAGCAGAATACCGGCACCGTCACCGTTCCCATCAGATGAGACGGCACCACGATGTGTCATATTCACTAAAAGATATCTAGCGTCAGTAACAATCTTGTGAGACTGTTCACCATGCTTATTTGCTACGAAACCGACACCACAAGCGTCATGTTCATAATCAGGGTCGTAAAGTCCTCGTTTGTCCGGAATCACATTTGCCCAAGATTTATGAAGATGGTGTTCATC tpg|BK006938.2|:154077-156022 7X251= 219=7X 
 tpg|BK006946.2| 235802 + tpg|BK006946.2| 236104 - INS GCCTGTGTTTGATCTTATGCAATAAGAATATATACAATTTATGTAGTAAAATACCTTTTCTTCTGCGAGTTGCAAGAAATAGAAAAGACTCCGATTGCGCATCGCCAGAATAAAATTTCACAACCACACTTTTTGGCTGAACTTTTTATTACCTGATTAAACAGAGAGAGAAAAGGTAGAGGTCAAAATTTTTTAAGCAAAACTAAAAAAGATGCAAAATCACGTGCTGAAAATCTAACATAAGGGTTAAGATTAGAGTTTTATAGGACTTGTTTTGTAATATTTCAAATACGAGCTAACCCTACTGATTTCAATTAGGTCTAATTTAGGGTTGAGCTGCACTGAAATTTCGGAAATTTTGGGTTATTTTAAATGAGACAGAAGAACTACAGAGATACGTTCTTCAGACTTTAAAGCTTATCTCCACAAAGAATTGGTCAAGAAATCATCCTAGAAAAACACGTTTGCTCACTCGATCTTAATCACATAGAGTGCTGGAACGGGAAGAAATGGGTATGTGCCTCGGTTTTTCTCATTAACCCCTTTTGATC tpg|BK006946.2|:234686-237220 7X5=151S 8S526=7X 
 tpg|BK006946.2| 790938 + tpg|BK006946.2| 790577 - INS ATCTTTGCCACCTTTAGGAATTCTGAAATCTTGAAGATAAATAAATGCTTTTTGGAGGCTTTGTAATCAGCACAGAATTTTTCTGGAGCCAAATTGAAAACAGTAGACGTTTCTTGGTTGGACTCCCAAGCATTATTTATGTATTCGAAGCACTTTGTAATCCAATTATCCGAATCATGTTCAATAACAGATTTGAATAATTTTTTCCACCTACGCCTTTTTTCTTCTGGAGACATTTCTAAACTTCTCTTGATACTTTGTGCTACATGATTTATATCCCATGGGTTTATTAAGATGGCACCTTCCTTTAGGACAGAAGAACTACCAGTGAATTC tpg|BK006946.2|:789893-791622 7X417= 315=7X 
 tpg|BK006946.2| 718822 + tpg|BK006946.2| 718895 - INS TTACCGTTAGCTTACTGCTTTCCGCTTGACTAATATGGGTTATTCTTGATTCATTATCAACATGTGATTGGGTAATGTCTGGAGATCCAGTTCTTACTTCTCTATTACTAGACCGGAAGGAATCTAGCCCATTACCATTGAATGCGAAATTTGTCTCATCATTTTCTTTAGGGGGAGTCGGCCTAACACTGTTAGCACGCTTAACC tpg|BK006946.2|:718396-719321 7X189= 194=7X 
 tpg|BK006938.2| 1172691 + tpg|BK006938.2| 1173303 - INS GACCTGGGACGTTATCTCGAAATGGATAGGCTCCCCGAGTTAAATTGTACGTTATCTCGAGTTACCATTAAATCGGTTATCAAAGCGGTCGAGGAATTTTCTGAGGAAACATTTGTAAAATTCATATCGTCTGTCACCAAAGTACAGTTAACAGC tpg|BK006938.2|:1172367-1173627 7X10=67S 71S7=7X 
 tpg|BK006938.2| 99672 + tpg|BK006938.2| 99375 - INS CTTTATTGTTAAGACGATTGCTGATATTGGCTGTGGATTCGGTGGGTTGATGATAGATTTATCACCAGCCTTCCCTGAAGATCTTATCTTAGGGATGGAAATTCGTGTGCAGGTTACAAATTACGTGGAGGATAGAATTATTGCCTTAAGGAACAATAC tpg|BK006938.2|:99043-100004 16S175= 140=7X 
 tpg|BK006938.2| 1196313 + tpg|BK006938.2| 1195868 - INS GAATATAGGCATCGCGAGGAATATAGGCACGGAAAGAGAAACTCGTATAAAGTGACCACGGATATCGAGAATTTGATAATTTACCCTTAACTGAAGTTATGGCACAATATCTGTATAAATTTTAATACATAATTTGCGGCAGGAATAACTGCAACAATACTCAAAG tpg|BK006938.2|:1195522-1196659 7X237= 146=7X 
 tpg|BK006938.2| 360842 + tpg|BK006938.2| 361127 - INS AAAATTTTTATTTACGCTTGTAAAATAATATTTTCATTTCTTCTATTTTCCTCTTTTCTTCGTTTTCTTGACTTCATACTTCATTTTTTGTTTGACTCCTTTTTGCGTTATGAAACGTGATGCTTCGATATTCTCATTGGTTTCTTAAAACTTTAGCAATATCGGACAAACAGCCGTATTTTTTATTCTTATTTTTACTGCTTGATACAGTACCCCAGTCAGTGGCTGTTGAAACTCTGCCACTTGCCGTTTCTGATAGTACTTGCTTATAAGTTTTCATTGAATGACTTTTTTCACCAGCGGTATAGCTCTGAAATAATT tpg|BK006938.2|:360186-361783 7X218=22S 1S1=236S 
 tpg|BK006938.2| 910999 + tpg|BK006938.2| 911513 - INS GTTATGGGTGGTATCTATAAAGGCTTCCAATTGAATTTCAAGGTTTTTGGCTCAGAAAGTAATAATACTGACTACGACGTTTGGGAAAGTTTTAAATTGGATGACATAGCTGAATTTCAACCATTAAAGTTTGTCTCTAGAAATGTTAT tpg|BK006938.2|:910687-911825 7X4=70S 66S6=1X2=7X 
 tpg|BK006938.2| 730119 + tpg|BK006938.2| 730401 - INS ATTTATCACCACTTCCATCTTCAATGTTGCATGCAAGTGTTCTCAATTTTGAATGGGAACCGCTCGAAAAAAATATTTCGGCAATTCATGATAGAGATTCTTTGATTGACATTATACTTAAAAGATTCATTATAGATTCAATGACAAATGCTATTGAAGACGAAGAAGAAAATAATCTTGAAAAAGGGTTACTAAATTCGTGGATAGGTCTCGATTTTGTGTATAACTCAAGATTTAATAGATCTAATCCAGCTAGCTGGGGAAATACCTTTTTCGAGTTATTTTCCACCATCATTGAT tpg|BK006938.2|:729507-731013 7X189= 53=1X96=7X 
 tpg|BK006938.2| 732531 + tpg|BK006938.2| 733021 - INS CCGCCAAGATCGATGGCTTTAAAGAATTCCAAAACTTCAGAATATCTAAGGAGAAGATACCGCCACCCGCTTTTGACGAAACTTTTAAAAAGTTTACGTTCATCAAGATGGGGAATAAATTGATTAATAATGTTTGGAAAATACCTACTGGTCTAGATAAAATTGAGCAAGAAGTAAAGAAGCCTGAAGGTGTCTATGAAGCAGCCCAAGCGAAATGGGAATCAAAAATTTCTTCTGAAACTTCCGGTGGAGAAGCGAAAGATATGT tpg|BK006938.2|:731983-733569 7X133= 179=7X 
 tpg|BK006946.2| 234712 + tpg|BK006946.2| 235198 - INS TTCTCAAAATGACGGTTAGCTGTGCTCTCATCTCCGACTTCTCTCTTCAATAAAGTACTGTAGACACCGTAAAGTACAGCACCTGCAAGTGCCAACAAGTTGCCTATCAGAACTTGCACGGCATCGTTATCATCACCACTAACGTCCGCGATATGGCGTTGGTAGCGCTGATGAGAATCTGATTTGGTGACCATGATTATGCCTACAAAGGAAATGAACGACCCGAGTACTTTGGACTTGCTCAACGATTCAACATGACAAATAGCACCTATGAACAAGGTGAAAAAGGAAGAAGTAGTGGAGAGGATTGTCTGCGATGCCACCGATGTGAATGCCAGCGAGGCATTGGTCACAAGGTTAGCTGTGAACCAAAGTATGCAGAACTCAGCACTTAACTTGATTGTTTCATATAACGTTAGCCTCTTCTTTTGGTTGGCATGCGTGCCTGCTTCAAGGTTTGTAAGCAGTGGGCTAGTCATATC tpg|BK006946.2|:233734-236176 7X6=134S 10S457=7X 
 tpg|BK006938.2| 861877 + tpg|BK006938.2| 862392 - INS TGTCTCTTATTCTTAGGAACAGCGTATCGTTATAAAACTCTCCTCGAAGAAATTTCCAATAAATACAGCATATCCAATTTTAAAAAATCTCTGGACTTCTTTCGTTTAGCTTCGTTGGTGTTACCAAGTGCTGGTGAGACGTATTCGCAAGCAGGAGCG tpg|BK006938.2|:861545-862724 7X77=42S 3S1=37S 
 tpg|BK006938.2| 339848 + tpg|BK006938.2| 340455 - INS TTCATCATCATGGAACTCCTTGTACTTGTGACTAGAATTTTTTATTATATCGCCAATATTTAATGATAAACATAATATAGTAATACCAAAAATAATTATGATAACTTATACAAAAGAAGTGGAAAGAAAAGGAAAGAAGTAATCAAAGTAACTCAAAAAAGGTTAATGATTACGATGTTACAATCGCTCTTGACTTATCTGTACTTGTGGAAACCAATGTCGTTAGCCTTTTCTCTGAAACATTGACGACAGATGTTTAAGTCGTACTTTCTGACCAAACCAGTGTGGGAGGAGCAGACACGACATTGACGGGAACCTTTACCGAATCTTCTTGGGTGGGAGAACCAAACGTTTTCGTGAGCCATTTTGTATATATTCTATAACC tpg|BK006938.2|:339064-341239 7X267= 361=7X 
 tpg|BK006938.2| 659103 + tpg|BK006938.2| 659722 - INS TTATCCTATACAAGGATAACGATGCCAACTTGAGAATGACTACACTCGAAGCTTCAGTACTCAAATGCACCTTAAATAAACAACATTGCGCCGATTTATCAGATCTTTACATTGTTCAGAATATAAATTCTGACGAAAGCACAACTGTACAGAAATGGATATCAGGTATATTGAATCAGGATTTTGTATTCAATGAGGACAATATCACTTCGACCCTGCCTATTCTTCCCAGTATAAAGAACTTTTCAAAAGATGTTGGTAATGGTAGGCACGAGACGAGTACCTTTCTAG tpg|BK006938.2|:658507-660318 7X11=250S 4S209=1X59=7X 
 tpg|BK006938.2| 1306915 + tpg|BK006938.2| 1307214 - INS AGTAGCATTGTACGTACTACATCAATTGATAGTTTTAGTATGAGTGAAGTAGAGCTTTCCACATATTATGACTTAAGTGCTGGCAACTATCCTGACCAAGAACTGATTGTCGATCGCCCGGCCACTTCTTCCACTGCCGAAACATCTTCAGAGGCAAGTCAAGGTGTAAGCCGTGAATCTAACACTTTCGCAGTATCTTCGATTTCCACGACAAACTTTATAGTTAGCAGTGCTTCGGATACTGTTGTTTCAACTTCAAGCACCAATAC tpg|BK006938.2|:1306363-1307766 7X173= 253=7X 
 tpg|BK006938.2| 1293017 + tpg|BK006938.2| 1293054 - INS CGTCTCTGCCTGAATCTGTGCCACTGGTTTGAGACAATGTTGCAGGGGCCGTACCCAATCGTTGACCTCTTCCACTAAAAGTTCTCGTTTCTCTTTGCGAAGATGGCACATTGGCAAAGTTGTTGTTGAATGTTGCAGTTTCATTGTGGGCACCCGTTATGCGAGCATATAGACTAGTAAACCACCATGGCGTTGAGAATTTCCCATTGGGCGAGATTCCGTAGGTTGGATCAGCTTTTCTGGATATCATCCCCCATATTGGCCCCAGTGTATGGGTATCTAAG tpg|BK006938.2|:1292435-1293636 10S167=43S 67S4=7X 
 tpg|BK006946.2| 363977 + tpg|BK006946.2| 364680 - INS ACCTTGAATGAGGCAGGATTGTTTTGATTTGCAACTTGATTGTTTCCAAATAATCCGCCTCCAACAGTGTTTGATGGTTTTGAACCAAACAGGCCACCCGAAGCAGGTTGCTGTTTATTTTGGAACAAACCTCCTGATTGCTGCTGCAAATTATTTCCACTTATACCGTTACTTTGATTTGTTGTGCTGTTAGAGAATAAGCTTGTATTTCCAAAACCAGTTGGTTTCGCTCCAAAAAGACTATTATTCTGTTGTGGTTGTTGTAACCCATTTTGGCCAAATGGCTGATTATTATTTTGATTGGTCTGGCCAAACAATCCACCAGGTTGGGACTGCGACTGGTTGTTTTGT tpg|BK006946.2|:363261-365396 7X448= 330=7X 
 tpg|BK006938.2| 1006071 + tpg|BK006938.2| 1006672 - INS CCTTGAGAGGAACCATGGATACACTAGTTTGTGTTTCCACTACTTGTGCATACACATTTTCTGTGTTTTCTTTAGTTCACAATATGTTCCATCCCTCAAGTACTGGCAAACTCCCAAGGATCGTTTTCGACACATCAATCATGATCATTTCATATATTTCCATCGGGAAATATTTGGAAACTTTAGCTAAATCACAAACATCAACCGCACTTTCTAAATTAATTCAGCTCACTCCATCGG tpg|BK006938.2|:1005577-1007166 7X133= 120=7X 
 tpg|BK006938.2| 422242 + tpg|BK006938.2| 422516 - INS CCGTAAATAGAAAACATTACAATTCTATGCTCTGTTGAACAAACGGTGTGATGATTTCTGGTGTTTCTGCTTTTATAGTACTGTATATTACGTTCCAAAACGTGGAGCTGCCTTTCTATGGTGTCTATAGAATTTTCCACACTGTCTTGCAAGGGATCGGTTTTAGAGTCTCTCAGGTTTCTCTGCGC tpg|BK006938.2|:421852-422906 7X3=91S 90S4=7X 
 tpg|BK006938.2| 1190012 + tpg|BK006938.2| 1190536 - INS AAAAGCTGATTTATTCAACGAAATGTTGACTTCAGCCGATGAGCCTGATCTTGAAAATGAAGCTATTCAAGAATTGTATGGCGACTTAAAATCAGCGCAGCCGAAATTCAAAAAGCTTATTGAGGAAGAACGCGATGACGATGCGCTTGTTAGTAATCT tpg|BK006938.2|:1189680-1190868 7X76=43S 14S1=168S 
 tpg|BK006938.2| 456357 + tpg|BK006938.2| 456355 - INS CCCCAATCTGTAAATGGCAGAGAAGTAAATATAATATTGTCATAAAGGTACATAGTTGAAAAGGGTATTTTTTTAAAAATAGAAACTTACAATAGTAGACATAAAGGGACTGTTTTTAACGATTATAGGTGTAAGACAAGGAAAATTCACAAATTAAAGTTTAAAACTACTGTAGGGATTCTTCTTGATCCGATTTATCATCTATTACATTCTCATCATAAGTGAAATCGTATTCTCCTTCGTATTCATTTGAGCCATCATCTATTATAAGCTTTCCCTGAGGTTTTTTTGCCAAGGCATCTTCCACTTCGCCTGTACTCGAATTTAGACGCGAGCAAATCAAGTAAAGGTAAGCCACTCTTTTCCTTTTCCTGTTGTAAAGAAAACCTATAAG tpg|BK006938.2|:455553-457159 7X315=4S 11S167=1X203=7X 
 tpg|BK006938.2| 269083 + tpg|BK006938.2| 269419 - INS CGTATAACAAGTTACAAATATATCCGCCCCCTTCAAGAGATGAATTGAGGAAAAGGTTCATTGCTGCTAGCGAATACGCCTTAGATTTTATGTGTGGAATGCTAACGATGAACCCAAAAAAGAGGTGGACCGCTGTTCAGTGTTTAGAAAGTGATTATTTCAAAGAATTACCACCA tpg|BK006938.2|:268717-269785 7X4=84S 81S7=7X 
 tpg|BK006946.2| 304326 + tpg|BK006946.2| 305009 - INS TTGTTGCTGTTGATCTGGTGGTGATTGCAGAACCATTCGGTAACGCAGTTGCAGTAGCGTTGGAAGGAACACCTACAGACGTGGAAGGTGGATTGGAAGCATTTGAGTCAGAACCGCTACTCTGAAAGGATTCTTGAACTTGATACATCTGAGGCTGGGATTGCAGTTGCTGTTGAGACTGGGATTGCGGCTGCTGATAATATTGCGGGTACGGCCACTGTTCAGGAACTACGTATTGGTAGGATACGGGCATCAGAGGTTGAACGCTCTGGCCGAGATATTGT tpg|BK006946.2|:303744-305591 7X169= 267=7X 
 tpg|BK006946.2| 238788 + tpg|BK006946.2| 239028 - INS CATGTACTTCTTAAAGAAGTTTTATGAAGTTTCGTAAGTATTGGGGGGGTTGAAAATAATCTCTCACGTTATACGCAATAAAAAATTAAAATTAAGGAGAACCAATCTATAGAAACGAACCATTGAATTTAGCTATATGACTATATACCATTACGTAATTTATATAAACAGCTTAATATAGCGAAAGCAAAGTAGAACGAAATTTCGGAGAGTTCTAGATTGTATAGAGCGAATGAGCATTCAATACACACGCGAAGGCAGTAGG tpg|BK006946.2|:238244-239572 189S54= 133=7X 
 tpg|BK006938.2| 1330734 + tpg|BK006938.2| 1331191 - INS AAGTTAACCATTTATGGAATTCTCAGGAGCAACGGGTCCCTTGGTCTTTACAAGTTCTTCCATATAATGAGACTATTGAGCAGATGGAAAGTGAAGGCAACCAGTTTCATGTCGTTACTTTGAAGTTAGACGAATTTATTGGTTACTCATCAGCTTACGAC tpg|BK006938.2|:1330398-1331527 7X15=1X43=21S 5S1=221S 
 tpg|BK006946.2| 495582 + tpg|BK006946.2| 494971 - INS AAGGTCACCTGCATACTGTGTATTTAGTGTATTTTGCTATATCAATGGCCATTGAATTGGGACTTTCCCGTATTACAAAACTACTAGAGCATTTAGGCAATCCGCAAAACTCACTTAGAGTGCTGCACATTGCAGGGACAAATGGTAAAGGTTCAGTATGTACTTACCTATCTTCTGTGTTGCAACAAAAGTCCTACCAAATTGGAAAATTTACCACTCCACACTTGGTGCATGTTACTGATTCCATTACAATCAACAATAAGCCGATTCCGTTAGAGAGATACCAGAATATTAGATTACAACTAGAAGCTTTAAACAAGTCACACTCTTTAAAATGTACGGAATTCGAGCTATTAACATGTACCGCATTCAAATATTTTTATGATGTGCAGTGCCAATGGTGTGTCATAGAAGTAGGCCTTGGCGGAAGACTTGATGCGACCAATGTTATTCCAGGCGCAAATAAGGCATGTTGTGGTATTACTAAAATCAGTTTGGATCATGAAAGCTTTTTAGGTAACACCTTGTCTGAAATCTCTAAAGAGAAAGCAGGTATAATAACAGAAGGGGTACCC tpg|BK006946.2|:493807-496746 7X3=239S 9=1X548=7X 
 tpg|BK006938.2| 287331 + tpg|BK006938.2| 287795 - INS TGCAGTCTACTCTTTGGGGGCTCCATTATCAGCTTGCGTCATCTCTCTACCATGGGCGGTTATTTGCATTCTCATTCACACAATTATCCAGCTGGTTCGGAACAACAACAAAGCACTTTATATCCTCACATGGATGCCAATAACGATTGGTTGTTGGAACTTTACAACGCACCCGGCGAATCTTTAACAACATTCCAAAACCTAACCGATGGTACCAAGGTCAGACTATTCCACACTGTTACAAGATGTAGATTACACTCTCATGACCATAAGCCACCCGTTTCAGAAAGC tpg|BK006938.2|:286735-288391 7X276= 273=7X 
 tpg|BK006938.2| 1403587 + tpg|BK006938.2| 1403955 - INS GTATCGTAGCGCTGCATATATAATGCGTAAAATTTTCTCTTTTTAAAAGATGTTAGTACGTTGGGTTTGGCTTGTTCATTTTTATTATCCTTTATTTACTTGTAAAAAAACGAAAGTGACGAAGTTCATGCTAAGATTGAAGAAAATTATTTATCGTATACTTT tpg|BK006938.2|:1403245-1404297 7X5=77S 76S6=7X 
 tpg|BK006938.2| 1019175 + tpg|BK006938.2| 1019787 - INS GTGCGTGATTACCATGATAGTGGTTGCCTAAATCCGGATATAAAAGCTAGCTTCATAGAACTCGAAAACTACGAGACTACGAACGAATTACAGAATGCTGAAAGAGAATTACTGATGAAAAGTGCCATGAATGTAGGCCTAAATTCGAATGGCAGGGTTTCATTGCCAGTGAAAAAAGTTACCAAAAAAATAGTTCAAAAT tpg|BK006938.2|:1018759-1020203 22S29=56S 95S6=7X 
 tpg|BK006938.2| 1446352 + tpg|BK006938.2| 1446527 - INS CTATAATATTGTACTTGCACTTAATTTTTGCAAATTATTTAATAATGCATCTTGCAAAACTTCCAGGTCCTGCAAAAATGTCACGACCATAATCTTTAATGGCTTTATAGTTTGTTATGCGCCTTGGCAGCGTGATCCGATCTTACTTGTTAACTGTATATCAGGTATTTCTGTTGGCATTTTTACAACTGCGAATGTATTTTTCATTATTTAGTAACAATTCTATTTACCCGGACAGCGTGTGCAGGTGATTTATTGATAAAGTCACTGGTAAAGACGTGCT tpg|BK006938.2|:1445772-1447107 21S127= 62=87S 
 tpg|BK006938.2| 671596 + tpg|BK006938.2| 671830 - INS CCTCTTTATTCTTACTCCCAAGAAGAATTCGAAAAATGCCAGGCGTTAGCTAAGAAACTAAAGAAGCAGTTGTTTGTTGAGAGTATCTTACTAGCACTCTGGAAGGATTCTTTTATTTACGACGAAAATTCAGTCATACAGTTACACCAACCAGTAATGTCATCGCTTGAAGAAATTC tpg|BK006938.2|:671226-672200 22S74= 63=33S 
 tpg|BK006938.2| 35847 + tpg|BK006938.2| 35867 - INS TGGACTAGGAGGCCTAAATTGGATGCAGTATATTTGTGAGAGAGAAATTTCGAAAGCTTGACCTAAAGAAGTATTGACCAGGTTACTAAAGTTTATTGAATTTTCAATAACAAATGGTGTAGAAG tpg|BK006938.2|:35583-36131 7X4=58S 58S5=7X 
 tpg|BK006938.2| 676896 + tpg|BK006938.2| 677645 - INS TGCATATAAAGTATTCAAAAAGGTGTTGAAAGCTCTTCCTGTATATGACCCTGTATTTAATGTACGCGGTTAAAAAATTTTTATATTTTTAAATAAGTATCAACTTGGATAATATGATCTTGCCCGCAAGG tpg|BK006938.2|:676620-677921 7X60=38S 4S1=211S 
 tpg|BK006938.2| 685052 + tpg|BK006938.2| 685123 - INS TTAAAGTTGGTTTGTTTTATAGTGGAAGTACGAAAGCTATATTCCTCATTATTCGTTTGTTTTTGGAATGTTTGTAGCAACTTCTTTCTTTCGGAATTCTTCAAATTACTTAAAGCTTTTATGTGAGGCTCCTTCTTAAACATAGCTGTACTAATCCTGCGCTACACTAATCTAT tpg|BK006938.2|:684688-685487 7X6=81S 83S5=7X 
 tpg|BK006938.2| 230056 + tpg|BK006938.2| 230202 - INS ATTCGACTAAACATACAAGGAAAGTCATTTTTTCTGCAACGTTTTTTTACCCTTTATGTATATATATTTACATATAAAATAAACCTCTAATCAATCAGTATTTAAAAATCGGAAGTAATGTCCATACGAAAGGGCTACGAGAATTTAACCATCTCGTTCTTTGCTAG tpg|BK006938.2|:229708-230550 7X33=50S 1S1=250S 
 tpg|BK006938.2| 378865 + tpg|BK006938.2| 379029 - INS TTCTCCGAGCGCAGCTTTAGTGTGCCCAAGTGGATCTGTTGTGTTGGTTTCCCTCAAGGAATCCGGCTGTGCTACTTTTATCTTCTTATGTGAAGGTTCATCATTATTTATAATGTCATCGGGTTGTTTTCTGATCGCGTCTTTATCTTGTGTGGGGCTTACTGTATTTGAAACCTTATTTT tpg|BK006938.2|:378487-379407 7X5=86S 85S6=7X 
 tpg|BK006938.2| 178576 + tpg|BK006938.2| 179017 - INS GGTGAATACAATGCTTTTGAAGATGTGATACATGGCATAAGGTATATCGACATAAGGGATCGGATGGTACTGGATGAAAATACTATATCGGCTTTGCATATTTTTCCAACAGCTCATAAACTGGGCCATGATAAGATGATGAGAAATGGTTTCTTTAGTGTATTTGAACTATTCAATCAAGTGTCTTCGGACTACGCCAGGAGAATTTTGAAGTCTTGGCTTATTAACCCATTAACCAATAAAAAACGGATAGAAACAAGATACAGCATCATAAGAACCTTATTGGATAAACAAAACGCCATCATTTTTAGTGACCTTAGCCAATCAATAAAAAGATGTCC tpg|BK006938.2|:177880-179713 7X13=16S 320=7X 
 tpg|BK006946.2| 738511 + tpg|BK006946.2| 739094 - INS TAAATCTAAAAGGAAGAAGAAAAAGAATGATAGTCCTGATTCCAACAGCATTTCCGTCCGCAAAGTTCTGTTGTCAGCTCCTTTACAAAAGTTTCTAGGATCTGAAGAACTGCCACGAACGCAAGTAGTGAAGATGATATGGCAGTATATCAAAGAGCATGATC tpg|BK006946.2|:738169-739436 5S2X11=71S 77S5=7X 
 tpg|BK006946.2| 134040 + tpg|BK006946.2| 134271 - INS ACTTTGATGACCTTGTTAGTTAACAATCTCGGCGGTGTTTCTAATTTTGTTATTAGTTCTATCACTTCCAAAACTACGGATTTCTTAAAGGAAAATTACAACATAACCCCGGTTCAAACAATTGCTGGCACATTGATGACCTCCTTCAATGGTAATGGGTTCAGTATCACATTACTAAACGCCACTAAGGCTACAAAGGCTTTGCAATCTGATTTTGAGGAGATCAAATCAGTACTAGAC tpg|BK006946.2|:133546-134765 7X4=342S 225=7X 
 tpg|BK006938.2| 268143 + tpg|BK006938.2| 268143 - INS GAATGATTATTTCAAAGAATTACCACCACCAAGTGACCCGTCGTCAATAAAAATACGTAACTGATATGATTTTATAAAATTTGTAGAATCTGTGTTATTGACATTAGATGTATCCTCAACATATACAAATAAACTTCTTGATCCGTCTTGTTTTTTGGTGTTGAATTTTAACTCTTTTCCATCATTATGGAATTCGTTTTTAGATTTTAACAACAACAATAT tpg|BK006938.2|:267685-268601 7X7=104S 106S5=7X 
 tpg|BK006938.2| 859931 + tpg|BK006938.2| 860310 - INS GGTGTATTGTCTGTACAACTTTTATATTCCTTTCGGTCCAAATCATTGGGCTTATTATCTGATTCGTTGCATATGGCCTTAGATTGCACATCTTTGCTCTTAGGTCTAATTGCTGGTGTATTGACCAAGAAACCAGCAAGTGATAAATTCCCTTTCGGTCTAAATTATCTTGGTACCTTGGCAGGTTTCACCAATGGTGTTCTGTTACTCGGCATAGTGTGCGGT tpg|BK006938.2|:859467-860774 7X246= 21=1X189=7X 
 tpg|BK006946.2| 720411 + tpg|BK006946.2| 721035 - INS GTGTACGAGATTCGGAATACACTCATGTTCATGACCCCATATCACCATATCCAGGAAATCTGGCAAGAACTGTTCAGGTAAAAATGCAGTATTCGTGTGACCTGTATGATTTTGATGGACGCACATTAAATTAAACCATTCACCTTCTCGCATAGTCGGTACTTCAAAA tpg|BK006946.2|:720059-721387 7X5=79S 75S10=7X 
 tpg|BK006946.2| 299014 + tpg|BK006946.2| 299437 - INS GCAATTACGAAGCTGCCAAGTTGTGAAAAGTTAAACGCACTAATTGGTCAAAGTAAAATCGTTCAAAATCTAACCGAATCATTCGATTTGAGTATTTGTCTCATATTTGGATTTGATGTAAGCGCTATGAAAGCAAAGAAGTATGGAGCAAGGGAGAAGACGGCCAATGCTAATCAGACGCACTCCAACATTGACTATGACACCGATGACGGCAATGAAAAGAATGCCATCGATAGCAAATCTAATGCGATCGGCGCACAAACTCAAAGCAATAAAGAAACAACGTCCGACAATGAGGATCTATTGATAAAGGAATACGAGGGAATGCTAGGCAGTTCAGGAGATGAAGGGGAAGGCGGCGGATACTTGAACCCTAATATCAATTACAATGAAGTAACAGATGAAGAACCT tpg|BK006946.2|:298178-300273 7X194= 206=7X 
 tpg|BK006938.2| 302290 + tpg|BK006938.2| 302833 - INS GTATAAAGAGGAAAATTCCACTGAAGTTGGTAAGCCCGGACCACAGCAGAAGCTATCGAAATCTTACACTGCGGTATTCAAGAAATGGTTTGTCAGAGGTTTAAAGTTAACCTTTTACACGACGTTGGCCGGCACATTGTATGTGTCATACGAGCTGTACAAAGAATCGAACCCACCCAAACAGGTTCCCCAATCGACCGCTTTTGCTAATGGTTTGAAAAAGAAGGAGCTGGTTATTTTGGGTACAGGCTGGGGCGCCATATCTC tpg|BK006938.2|:301744-303379 21S87=32S 128S5=7X 
 tpg|BK006946.2| 684337 + tpg|BK006946.2| 684243 - INS GCCTTGTCCTATTTAGCCCTATATCTACGTATAGAAAACTGTCAATATGTCATTACCGTTCTTAACTTCTGCACCGGGAAAGGTTATTATTTTTGGTGAACACTCTGCTGTGTACAACAAGCCTGCCGTCGCTGCTAGTGTGTCTGCGTTGAGAACCTACCTGCTAATAAGCGAGTCATCTGCACCAGATACTATTGAATTGGACTTCCCGGACATTAGCTTTAATCATAAGTGGTCCATCAA tpg|BK006946.2|:683743-684837 7X8=1X49=1X178= 4S224=7X 
 tpg|BK006938.2| 912402 + tpg|BK006938.2| 912429 - INS CAATGGATGGTACGGATAAGGGAGTGAAAAATCCAAGACCACTCGAAAAAAAATATAGTAGCAGTTGTTTTGAGGACCGTACGCCCCTTAACTTGGATGATGGTCATTTCAGTGAATGCAATCATTTTTCTACATTAGATGTGTCTAGCTTTTTTCATCTCAACGAGCATGTGCATAAAATCGACGAAGTAGAGCTCGATGGACCTGATCGCACCTTTAGTCTAGACA tpg|BK006938.2|:911932-912899 7X146=25S 3S1=208S 
 tpg|BK006946.2| 349664 + tpg|BK006946.2| 349470 - INS GGCCTGGGATGATCAAAGTAGCATTGGCTTCTCTTTCAGCGTTTTGAATGTTTTCCTCGTGTGGAAGTAGAGTAGGTGGAGCAGGTTTCTTCTTCTTTGAACGTGGCTCCAAGTCATGACTCTCATTAGATGCTTTGGACTTATCTTCTCTCCTCTTCTTTGGGCTGTTCTTGTCCTTCCCGTTTTTATCCTTGTCGTTATTAGTACTGTCATTATTGTTATCATCTTCATATTCGTCGTCGGACAATAGTCTAACCATTTT tpg|BK006946.2|:348932-350202 7X151S 246=7X 
 tpg|BK006938.2| 923680 + tpg|BK006938.2| 923514 - INS TACTCGTGATCCATAATGAAAAGAGAGTATTACAAATAGACCTAGTGTTTTCAAGTACAGTTTTCTTAACTACTCCGAAAATTGTCCTGGTAATTCTTTGCAATGCAAAATTGAAAGAGAGACTTTTAAACTACTAAACCCTTAACAGTAGAACAACATTGTCTCATTAATTTTTGAAATTTCGCTTTCTTCCCATGCCTTAGGCCAAGTTCTCATCCAATGCGTCGAGTCCTTAAAAAAAATTCGCCCGGGTAAACTAAAACTT tpg|BK006938.2|:922970-924224 7X163= 133=7X 
 tpg|BK006938.2| 346321 + tpg|BK006938.2| 346441 - INS GCCTAAGCATCAAAATGCGTTGCCTAACTCAAGCGTATTAATGGTTGTGTTGCGACTTGCATTCTTTCATAATATCCCAAAAAAAGTTAGACCGGTTGCTCTTTTGACTGCCGCAAACATGGTTAGAAGTAATGAACATGCACAGCTAGAGTTTAGTAAGATCGATGTTCCATATTTCGATCCTTCATTACCT tpg|BK006938.2|:345921-346841 7X4=227S 97=7X 
 tpg|BK006938.2| 181375 + tpg|BK006938.2| 182098 - INS CCTTCAAAACTAGATGGCAATTCGCTGGCTTGCCTCCAAATCTTTTTTGTCGTTAAAATCTTTTCCATGACCGGATGTCCCTTCATAGATGTGAAATCTTCATTATTATGGAGTTCGTGCAACAAGATACTATAGTAACATGATATTGTGCCTAGGTAACTTCCAAGTGCAATTAGCTTTAATTTATTGAACTCATTTTCCTCAGATTTCTTTAATTCGTCAAACTTTGGAGCTAATTCTGTGAATTCTTTTGAAAGTGGAGCAAATTCAGGAAACATTGTCCTTAAATAGTTATCCCTTGCTTCGTCATCCATATTTAGAATATCCGTTATGGAAGTTTTAGTATCAGCCTGCTTGGTCGAGTTCTTAAATTCACCCATGTCAAATTCTTTGGCACTTTTGACCCACTCTTCTTCTTCTTCTTCATCTAAGT tpg|BK006938.2|:180495-182978 7X9=12S 217=7X 
 tpg|BK006938.2| 940467 + tpg|BK006938.2| 940755 - INS TGTTTATACTCGGAGACAAGAAGAGAGATATGTGTAGGAAGCTTTTGTCTGTTCACGTAATCATTATCCAGTGTTCCAC tpg|BK006938.2|:940295-940927 7X7=32S 37S3=7X 
 tpg|BK006938.2| 945761 + tpg|BK006938.2| 946446 - INS AGACAACACGGTACCAAAGTTATACAATGACTGTGCACGCAACGTGGAAGGAAAAAGTTCAATTAAAAAAAGATCAACTGAACAGTAAGATAAAAGACGAATGGAAATTAAACAGCACAACTATAACGAGGTTGAAG tpg|BK006938.2|:945473-946734 7X1=1X7=59S 63S6=7X 
 tpg|BK006938.2| 1312784 + tpg|BK006938.2| 1313551 - INS AGGCGATTGAACTGATTGGGATAGGGAGTTTTTAAACGATGAGTATGTTCTATATTATTCTAATAAAAAAGATGATACTAATCTAGCACAGAATCACATACCACCATTTCCACTAAGATTCTCATTCGCCCAAAGAGCAAAAATAGAGATCATTCGAATCCTATCCATAGCATATGAGACGATTTACTGTGAGAAGAATAAGAGGAAATTGGCAACGACAGATCAGAGACACAACCTCTCTGTCCTAAGTGTTTTTTCTCCCTTGATAGAGGGCTGGCTCAGTAACTACAG tpg|BK006938.2|:1312188-1314147 7X185= 4S269=7X 
 tpg|BK006946.2| 538200 + tpg|BK006946.2| 538218 - INS GACCTGAGTTCGAAGAGTAGTAATTATTGAATTCTAAACCTTTTTCCTTTCCATTTGAAGAGGAAAGCAATTCAGAAGTTTGATTCCAGTAATTTTTATTTTCTAAGTTATGAAAAGTTGTCGCCGCTGAACCTGTGCCAACATTTCCATCCCTTTGATTTAGCCAAACTGAATTAGCAGCAGCCGTGACCTCGTTGC tpg|BK006946.2|:537790-538628 7X10=89S 94S5=7X 
 tpg|BK006938.2| 144450 + tpg|BK006938.2| 145047 - INS AAGTAGAAGGACCTTGGGCTTAGCCTTTTCATTATCATCTACTAAAATATATGCTCTCCATATACTAGGACATCTTTCTTTTGAGTGTTTCTTACTCTTACAAAGAGTGCACTGAACTTTTTTCCATTTATGTGGACATTGTGACCTGTAATGACCCACCTCATCACACTTTGAACACTGGATAGCCTTCGGACAATGTCGAGAATAATGATCATCCGTCGCCCCACAGTACGAACATATTATATGGGGACAATCCTTCTTCAAATGACCTCTTTGAGAGCAATTATTACATTTAGGTGCTGCCTCTTTAATGGCATCCTTGTCATCATCGCTTACGCCAAAATATCTACCCTGCCCTCTAAGAGCTCTTAATTCGTTGGGATTACTATTTACTTCCTCTATAGAAGGTGCTACAAGTTTATCTGGAGGAGTTGTGGGTGCCGTATCGACGACAAATGGTGCCGTATTTTTTTCCATGACTGCGAGGAAGTGATGTAAGCTGCTATCGTTGTACAGGTAAGGTTTAATTCTCTCTGATGCTGCCAATAGTCATAACTTTTTTCGAAATGTTTCTTCCCATCCCATTAG tpg|BK006938.2|:143260-146237 7X229= 294=7X 
 tpg|BK006938.2| 150971 + tpg|BK006938.2| 150928 - INS CCCTCACAGGGTGCTGGACATACTCTTCCAGTGAATTCTGGGAAATTGTTTGTCTCTAGCAATTTGTCCAGTGCCAACTTCCATTGGTTCTTGAATAACAATTCATTAAACTTGGGGATAATGTTAGATAGGGGACAA tpg|BK006938.2|:150638-151261 7X2=67S 65S4=7X 
 tpg|BK006946.2| 156308 + tpg|BK006946.2| 156322 - INS TAAATCAGCCGATCCGCTCGACTTATCTACAGTTTTAAACTTACGAATAACGGCCTCTTTCAAATAATAAGGCAATTCATAAACGATGGATTTATTTAGTAAAACTTCGATATCCATGATCTCCTTTGTTAAACCTAAGTAGTCGTGAGCAGTTTGGAACGTAACATGGTATAGCTTGGTGAGAACCATCTGTATGATATGGGAAGCAGACCGTGGGTATTTTGCGGTTAATTTGGCAAACGATTGAGGTGGGAT tpg|BK006946.2|:155784-156846 7X100=27S 4S1=367S 
 tpg|BK006946.2| 398803 + tpg|BK006946.2| 398915 - INS ATTCACGGCATGCGCTACGGAATACAATCCTAGCCTGCTTGATGGCAAAAAAATTGCTCCATCACTGATAAAACACCCGGTGAGCCTAAAAACCATACTAGTTGATAGCAAATTAAAGTTTGATGGTATTAGGGGAGTGAATAAATGGTTGATGGAATTCGTTGCAAGACGACAA tpg|BK006946.2|:398439-399279 7X7=80S 83S5=7X 
 tpg|BK006938.2| 800154 + tpg|BK006938.2| 800499 - INS CCATTAGTCTTTCCTCATCGTCATTCAACTTATCCATATTTTCCAGAGTTAAAGGAGCCGGCGTTTCTGCATTTTCAGAAGCCTCGGAAAGTTCTATGGCGGATTGTTGTTGATGATTTTTTGTCGATAAGGATACTGCTGAAGAGGTACTTTGTTTGAGATCGATTTTATCATACACCGAACTAATAATTTGTGTCAAGGTCGCCTGTGCAATACCTTGATTGGAT tpg|BK006938.2|:799686-800967 7X186=19S 1=285S 
 tpg|BK006938.2| 1018134 + tpg|BK006938.2| 1018233 - INS TGTGACAAGTTGAAAAGTCCACCAATTTCACGTTGAATTAGGATTCATATATGAAATTCTAGTCATTAATTAGAATTGTAAGTTTCTGAGCTTTTTTTTCCTAGTAAATTAAACTTGTCTAATACATCCAGTTGTGATGTATTCTATATCTCAGTTCTACAGTAGCACGAAGTTTCCCGGCCTCTCTATTCAATAAATTCAGCTATCGCTGATTATCAACAGCAGCAACGAATAAAGCATAAAAGAACAGAAAAATTCTTCTACAAATTTATTCTGTAAAGATTCAGCTTCTTTCGTGAATTTCTAAGTTCATGAGGGGAATTTAAGTATGGCGTTTCTTCGTAGCGCCATTGTCTTGAGC tpg|BK006938.2|:1017398-1018969 7X322=16S 1=184S 
 tpg|BK006938.2| 348172 + tpg|BK006938.2| 348148 - INS TAGAGAATGAAGACTAATGAACATATTTCGAAGGAACTTGTTGAGTACAAATCCCGCTTTCAGAGTCATGACAATCTAGTAGCGAAACTAACAGAAAAATTGAAATCCTTAGCAAATAACTATAAGGATATGCAAGCTGAAAATGAGTCTCTAATAAAAGCTGTAGAAGAGTCAAAAAACGAAAGCAGCATACAATTGTCT tpg|BK006938.2|:347732-348588 25S82= 34=74S 
 tpg|BK006946.2| 38384 + tpg|BK006946.2| 38622 - INS CAAGTAGGATATGTTTTGACAAGTCAGCTTCTCCATATATGCCATTCCGAGTACTATACCAACAAATATTCATCATTTTTCTATGGATTGGATTGGTTCTGTTTTGGGCGTGATAGGTCTCATTTTATTAAATTTTGTGTGGAACCAAGCTCCTATATCGGGTTGGAACCAGGCTTACATCATCGTAATTTTAATCATTTCTGTGATTTTTCTTGTCGTTTTCATCATTTATGAGATTCGATTTGCCAAGACTCCACTATTGCCGCGCGCAGTTATAAAGGATCGTCATATGATTCAAATTATGCTGGCTTTATTCTTTGGATGGGGCTCTTTTGGCATCTTTACGTTTTATTATTTCCAATTTCAATTAAATATAAGGCAGTACACGGCATTATGGGC tpg|BK006946.2|:37572-39434 7X171= 5S370=7X 
 tpg|BK006938.2| 371372 + tpg|BK006938.2| 372123 - INS CTATATATATAATTCTTTTCCCAGTATTTTAGGCAGAATATAAAAGCTTTGAGGCTTTAAGTGAGACAAAAGTCTTACCATAGCAACACGAGGGCTCGCCGAAACTTCCATCTAAAATAAAGAGTGCCCATTAATGTCCGGAAAACCACCAGTTTATAGATTACCCCCTCTTCCCAGACTAAAAGTGAAGAAACCTATCATTAGGCAAGAAGCGAACAAATGTCTTGTTTTAATGTCAAACTTATTAC tpg|BK006938.2|:370862-372633 7X172= 233=7X 
 tpg|BK006938.2| 380405 + tpg|BK006938.2| 380501 - INS GGAAATGTTGAGGCAAAACATTTGGGTGGTTCGCATCTTGGATAAAATTGTTCAAGTTTTCCATACAAAGCCTTCTTCAATTTATTGTCACCTTGGATTCCCAAGGATACTTCCAGTAATTTGTAGTACTTAAAATTATCTGGATTTCTCTTGATCAGAGTTCTATAAACAATGGACGCGTCTTTCAATTGACCCAATTTCATGTAAATAGTTGCTTTTCTCTCTAATAAACCAAATTTATCAAAGACGCATGGCTCGATATCATTCAAATGTTTCAATACATTTTGTAACTTGTCTTGGTTATCACTGGCAGCTTTATACATAATGTCGTTTTTGTACATTAAACACTCGCTGTGTTCATATTTCTCGGAATCAGATATTTTTCCCTCAGCGAGTTTTTCAAACTGAGATAAAGTGTTAATAGCTTGTTGCCTCTCACCGTTCACATCTTGTGCCACAGCCAATGATGTCCAGTTGGCACGGTAACCAAGGAATGCTTCCCAATATTTTTTCCTGGACACTAAAGCATTTTTGAAATCGCCAATTTGTGATTGCAAAGTTGCTAAGTCTCTATATATTTGCTTGTTAGTGGAC tpg|BK006938.2|:379203-381703 7X6=152S 1S575=7X 
 tpg|BK006938.2| 788646 + tpg|BK006938.2| 787955 - INS CCCTTAACATACTTTGATCCTTGCCCGTATCACTTATTATTTGGAATAATTGATTGATTTTCAAATAATACGACAGCTCCACGCACCCTTGACTTTTATCTTGATTAGTATTGTTTTGTAATATAAGCCTTTGAGAATGAATGATTTTACTAATCATATGGCCAGACAACTCGTTCAGTTCATTCTGAAAGCCATTCATTTTGATGGACATCCATCTTAGGATTGGATTTTCATTGGATGATGAAGTTGTGTTCTTGTTACCACTTTCACTTTCTCTTTGATTATTATTGATAAAGTTTTCTAAGTTCAACAATTTTGAAAAGAGGGACAAAATTGTTTCTTGGGGTTGGTCAATGTTAAAATTTGAATTTATTAAACTGTTCCAAATCAGATCTTTATACGTGACTAATAAATTTTCTATTTGAGTCCAAATTCTTTTTATAACAAGAGATTGTGAAGCATCTGAACTCTGGTTGAAACGGCGACGGAGCGTAAGAC tpg|BK006938.2|:786945-789656 7X3=198S 1S482=7X 
 tpg|BK006946.2| 795185 + tpg|BK006946.2| 795794 - INS CTCATCTTTTGGCCATGGAGGATTCGAGATTGCTCATCACTTTGATTCTTGTGTTTGGAGTTATATTTCTGAAAAAATTCTTCCAAAGTAATCAGCATCCCTCAGCACAACGCTTATCCGCTACAGGTGTAAACGCACACGGACGTCCTCAGGGCTCCACGCAGAATGCCTTGAGAAGGACTGGTAGAGTCAATGGAGGTCACCCCGTGACTACTCAGATGGTGGAAACAGTGCAAAATCTAGCCCCTAACTTACATCCTGAGCAAATTAGGTATAGTTTGGAAAACACAGGCTCAGTCGAGGAAACAGTGGAAAGGTACTTGCGTGGTGATGAATTCAGCTTTCCACCTGGGTTTGAG tpg|BK006946.2|:794453-796526 7X77= 180=7X 
 tpg|BK006938.2| 1080777 + tpg|BK006938.2| 1080885 - INS GGCCAGAACTGCCCCAACGTACGGACCAGCTTAACGGATATCTGGCGGTATGATTCTGGAATATTTGACCTGGTTGTTTTCTGAACCGTCATCAAGGAAGTCAAAAATTAACATGTTGTCGATGGTTTCATTCAGATTGTCTTCGTTAATGCCGTCCTGACCCAATGCCGGCAGTGTTTCGTTATGGGGAAACATCCACTCTCTCCATTGAGTGGTCACATTGTCGCAGAGGTCGTAGAGGATCATTTTTAGCAGGGTAATATGG tpg|BK006938.2|:1080233-1081429 7X175= 133=7X 
 tpg|BK006938.2| 1459603 + tpg|BK006938.2| 1459457 - INS ACCTACGGCAGGCGATTGTCGCCAATGGAAAGCTAGCCGATACTTTTTCCGTCAGCTTTGCGGGTTTTCTTTTTTGCGGCCTTGTAAACGGCTGTGGGAAAAGCGAAAAAAAGCAATGAGTTGGGAGAAATGGATGTGATTACATGAGCAACCAGTAGAAGATAGCATCAACCGCACACATGATTAGGATGTAGACGGCTATTACCTTGGACTTATTTTGTTCAAGTGCGGCTGTATGGACA tpg|BK006938.2|:1458959-1460101 7X5=144S 227=7X 
 tpg|BK006946.2| 43386 + tpg|BK006946.2| 43958 - INS TTATGACTAATTTCTATTATTGTCAGTGGAGTTTTTGAACAGATCACCTTGTGAATCTACAAACTGTCCTAAAGTATATTGGAGCAGGACATTGGGTGATGGCGAAAACTTTGGCACAAGGAAGGAAACCTGGAAGCGGCAGAAAGCCCGGAAAAGGGAAGACGTTGAGAGAGGGAAGAAAGCCTGGCAGTGGTAGGAGGAGGAGGCAAGATACTGGGGGTAAAGAGACCGACGGGTCTCAGCAAGATCAGGAGTCGCGTCTTATTAGTTCCAGGGACATGGAAGCTGTGGACGCACTGAGAGAGTTGACGCACAGCCCGTCGTCTCACTCAGCTCATAATTCATCAGCAGCACCACCGCCGCATGCAGCAGCGG tpg|BK006946.2|:42622-44722 7X267= 364=7X 
 tpg|BK006938.2| 1129519 + tpg|BK006938.2| 1130172 - INS AAAATAGATACATGTCAGGCAAACACAATGTATTCCAAGTTTTATTCTCCAAATATTCTGGCTGTAGGCTCTAGTGAAATGGATGAAAGCTCGTACTCGCATCACTCGGACGTAGAAATAGGGGTTGCTGTTATTGATAGATTCACCTATTACTGTTTGGATTTCCTAGAACAAATCGATAAAAATTCCACGTTAACTTTGCAGGACCTCTTCGATTCATTCACCTTCGAAAAGATTCACTC tpg|BK006938.2|:1129021-1130670 142S175= 121=7X 
 tpg|BK006938.2| 1416675 + tpg|BK006938.2| 1416569 - INS CGTGTAGGATCAGTAATTAAAAATACACACTATTCCTCGTTGTTATTTCTTAAAATTAGTTCAAGAAGAAGGGGTAACCCCTAAGCTTCTTAAGTTCACCACAAAAGTATTACTGGATAGTGAAACAACAACCACCCATAACATTAGTTTCCTAAACACTACGGCGGTATTCACCTAGACGCCATCCTAGAAGGCTACAAAGTGATGCACGTATGATGATATCGGACATTAGAGCGTATACATAC tpg|BK006938.2|:1416065-1417179 14S115= 123=7S 
 tpg|BK006938.2| 71396 + tpg|BK006938.2| 72064 - INS TAGTTTGCTGAGTTAAGGTTTCATTTCTTAACTTTCTTTTTAGGTTTTCTACAATCTCCAAAAGAGTAGTATCATTACGCTTAATGGTGATTTGAGATAAAAGGTTTTGATAATCAGAGCCTAAACGATTAACAAAATGGTTAATGAATATAGCACCAATATGAGCATATATAGCT tpg|BK006938.2|:71030-72430 7X6=82S 83S5=7X 
 tpg|BK006946.2| 221344 + tpg|BK006946.2| 221850 - INS TTAACAAGACAAGCGGTTAAAAGGCAGAGAATCGCCACTTCGAAGTCAACCACTATAATACAAACGGTATCTCCACCATCTCCGCCTCTGGACGTTCATGCTACGCCACTAGCATCCAGAGTCAAGGCGGACATACTTCGTGATGGAAGCTCATGTTCTCGTTCTTCCTCTTCTTCACCGCTGGAAAATACGCCGCCAAGGCCTCATC tpg|BK006946.2|:220914-222280 12S190= 7S6=7X 
 tpg|BK006946.2| 229072 + tpg|BK006946.2| 229158 - INS TATCCAAACTTTAGCTTTGGCCCTAGGTGTTGGTTTCGTTCCAGTCAGGAAGGCAGGTAAGCTACCTGGCGAATGTTTTAAGGCTACGTACGAAAAGGAGTACGGTTCTGATCTTTTTGAGATACAGAAAAACGCTATTCCAGCAGGTTCCAACGTTATCATTGTTGATGACATTATTGCCACTGGTGGTTCTGCTGCTGCAGCCGGCGAATTAGTTGAACAACTCGAAGCCAACCTTTTGGAATATAACTTTGTTATGGAGTTGGATTTCTTGAAAGGCAGGAGTAAGTTGAATGCTCCAGTGTTCACTTTACTGAACGCTCAAAAGGAAGCGTTGAAAAAATGATATGTTTCACGTCCTGACCCATATTCAAGCTTCCTTTCTGCCGGTTTCAAGCAATTTATTTTTCTTACTTCTCCTTACTC tpg|BK006946.2|:228206-230024 7X381= 213=7X 
 tpg|BK006938.2| 820274 + tpg|BK006938.2| 820583 - INS GCTTTTATGTTAAACGCGAAACTGCCGCCACTTCGCTTAAAAAAAACACTGGCTGAAAAAGAACGATGCAGTTTAGTAACTAAAGTTTTTTCTAGCTCAGGCTTAGAGTTCGATAACAACAAGTCACATTCGAGTGCTCCACTTATAGCAATTTTTCTTTTGTGTATTGGTTTGCTCCTGTGTGCTCAGGCTTTTCGTTTGTTGTGAGAGTATTGTTC tpg|BK006938.2|:819824-821033 7X9=100S 101S8=7X 
 tpg|BK006938.2| 721911 + tpg|BK006938.2| 722496 - INS TTTTTTATGGCGG tpg|BK006938.2|:721871-722536 7X5=1S 7=7X 
 tpg|BK006938.2| 692889 + tpg|BK006938.2| 693183 - INS TAAAAACCAGATTCGATCATCAGAGCTTAAAATTGTTATTCATAGCGGCACAATAGCAGAAGCCACAGAATATTACCTAGAGGTTTTAGGTGAAAGGAAGGATTTTTTTAATTATTTAATACTTTGAAATAGAAGTCAAGCCTTTCATTGCTTATTTATATCAGACC tpg|BK006938.2|:692541-693531 7X131=15S 2S1=191S 
 tpg|BK006938.2| 349331 + tpg|BK006938.2| 349997 - INS GATCAATACAAAATAACTAGAAATGACGAAAAGCTTCTATCAATAGAGCGAGATAATAAACGAGACCTGGAGAGCTTGAAAGAACAACTCCGGGCTGCACAAGAATCCAAAGCTAAAGTTGAAGAAGGGCTGAAAAAACTTGAGGAAGAATCTTCAAAAGAGAAAGCAGAGCTTGAAAAGTCTAAAGAAATGATGAAAAAGCTAGAGAGTACGATTGAGAGC tpg|BK006938.2|:348873-350455 166S90= 111=7X 
 tpg|BK006938.2| 365965 + tpg|BK006938.2| 366273 - INS GTGCTGTGCAACTTCTGGTAAAATCAAAAAAAGTAAAAAAAACGGCTCATGCCAGCGTGCTTCCTGTCAATAGCGGTTGTTGATTTTTTCGCTTCATGCCTAAAAAGAGAAACGAGACACAGAGAGAAAACAAGAATCTAGATTAATAACGTAGGGCAGCGTAACAATAATTTACGCAGAAATGATGTGTATTATTAGGGCATAAATAAATAAATGTATGTATGTGTGTGTATGTA tpg|BK006938.2|:365479-366759 7X297= 42=1X179=7X 
 tpg|BK006938.2| 973649 + tpg|BK006938.2| 973875 - INS GCATCTTCGTCTCTGCCAATGACAGGGTCTAATTTACCGTCGCGCGCTAATTTTGTCAAGTTTGTACCAAATTGTTCTAAAGCTGGCTTTTCCGGTTGCTGATTGGCATCCATCCTCATTTGGACGTACGTTCTTTTGAAATTGGGCAATCCATATGAGCTCTTGAGGGCGCAGGTTGAAATAGCGACTTCATTTAATGCATTTGTTTTTATATCTGATAGAAGTTTATTGGCTACTCGAGGTCTTGCATTAAAACTGCAAATAGATCTTTTACACTGTACAATAGTGTATATTCGTGGAGTACTTCGCCTTAATAGTTGCGTTCTCTGTAAATATTTTTGTATTGGTGCTTTTGTAGCT tpg|BK006938.2|:972915-974609 7X15= 180=7X 
 tpg|BK006938.2| 1254542 + tpg|BK006938.2| 1254549 - INS AATATCAGAATTAGTCGGTTCATTAACTAACTTTGTCCTTTTGTTACTGGGCGCCTCAGAAATCTCAGTATCAACTGGCCTCTTCTTTGAACCATTGATCGGTTCAGCATCGATGGTGATCTCACC tpg|BK006938.2|:1254276-1254815 7X5=58S 59S4=7X 
 tpg|BK006938.2| 715015 + tpg|BK006938.2| 715225 - INS GGGTTTCTCTACTCGCAGAAGAGGAGTGCTTTTTCACATGAAGGCCATCGGGAACAAGAAGAAAAGCCGTTCACGTAAGAAAATAGGACCCTATATCCGGTCAGGATCACTCAAGCTGTATGTAAATGTAATATAGACAAAGCACCTTTAACTGCTAAGAATTAATTATAGTGTCGGAAATATAACATAACTTGCTTACTTCC tpg|BK006938.2|:714595-715645 27S81= 29=80S 
 tpg|BK006938.2| 663865 + tpg|BK006938.2| 664109 - INS ATACCTAAGAAGTTTCCAGACTTGATTATTTTGATCAGCGTACCATTGTTTTGGAATACCACCTAGCAAAGTCACCTGTGAACATGCTGAAAGCTCTGTAGGTGAAACATACGACAGTCTAAACGCTGTGAAGGAATGCCGGGGAATGGTGAAGACCTTGACATTTGCATTTTGTGGTGAGCTGAAGCTAGTCACTC tpg|BK006938.2|:663457-664517 7X11=87S 94S5=7X 
 tpg|BK006938.2| 929206 + tpg|BK006938.2| 929219 - INS GGGTACAGAAGTATATTATTATTTCTCTTAATTATTTATTTATTTAACTAACACGATGAGCACTTTTAACTGCAATGGTTAAACTGTAGCAATGTTGGTAAAAAAGCAGGGAAAGTTCAAAAATAATTTATGTATTTTTCCTCGGGGGTACAGAAAGTAAAGAGAGAGAAACGTATGAGTATATATAGGCTAATGTAATATGTAGTGG tpg|BK006938.2|:928776-929649 7X258= 195=7X 
 tpg|BK006938.2| 582844 + tpg|BK006938.2| 582789 - INS CCTTCTAGTATGGATAATATGTATTTCAATCTAAGGGTTCTCAGGAATGGGAGATTGATTTCTCGTGGGTAAGATCCTCTATATAAATTTGGCTGTACAGTCGAAAATTGTAACGGAGTCACTAGTGTCATTTTGATACATATAGCTTATTCTAGATGTGTGAACTGGGTATTCAT tpg|BK006938.2|:582423-583210 7X11=77S 83S5=7X 
 tpg|BK006938.2| 1273039 + tpg|BK006938.2| 1272269 - INS CCCTTGGGTATTAAGAGGGCAAAGAGGCCCAGCGGGAGTTAATTTTTCTTCCCATTCAGGGTCAAGACTCCATCGAAACTGTTTCAACATTTCAGCCAAAGAAATTCTCATTTCTGTTAGGGCTAGTTTTTCCCCTAGGCATGCTCTTCGGCCTCCATGGAACCCAGTCACAGCACATCTGTTTTTCGCCATTCTCCAGTTTTTCCTTATGGTTTCGATATCTGAACCCCATCTTTCTGGTTTAAAATCATCTGCTGTTGTGCCCCAAGTTTTGGGAT tpg|BK006938.2|:1271699-1273609 191S12=28S 261=7X 
 tpg|BK006938.2| 753106 + tpg|BK006938.2| 753557 - INS GCTTCTCTACCATCTAGCAATCTATGATCATAAGTCAAAGCCAAGTACATCATTGGTCTTGAGACAATTTGTCCATTAACAGTGACAGGTCTCTCTTTGACACCATGCAAGCCTAGGACGGCTGTTTGTGGTGAATTGATGATAGGAGTACCGTATAATGAACCAAAAAC tpg|BK006938.2|:752752-753911 7X85= 155S6=1X2=7X 
 tpg|BK006938.2| 506715 + tpg|BK006938.2| 506280 - INS CGGTGTTAGTGCTCTTCTTGTTCCCATCTACGGGTTTCACGGAAAAACTACCCCGAAAAAGAAGCACAGCTTTATAAAAAGACCGTATTAATTTGCTTTATTGGGTAATAACGGGGCATTCGGGACATACAATCATACGCTAGATGCTGCGTGTAATAATTAACATTGTAAATCCCTATCTTTTTTTTTTATATAAGTAGAGTACTTTAAAAAGAGTGGACGACTGAGTTCATATACAAGCAGACGCCCTTTCATTTAATCTCAATCTTGTTTCAGGCCGGCTTTTGTCCATAACTGCTACGCTGCGTAAAAAAAAAATAAGAGAAATTGAAAAATATGGGCGTCGTCTAAGGATGGTAACTAGCTTCATTATAC tpg|BK006938.2|:505516-507479 7X4=208S 352=7X 
 tpg|BK006938.2| 957887 + tpg|BK006938.2| 958430 - INS TTTTCTGTCAATGATGGATTGTAATAATATTTCAGGATAAATTTCTCTATGAGCTGTAATCTTGATCTATTCTGCAAAAAAAACTCAAAGTTCAGACTCCCTAGTGAATCAGCATACGTGAAATATAATAAAAATATTACAGTCGTAAGGGGTTCAATAGACGCTAGTTTTTGCACTGTAGATCCAGAGACGTATAGGATTAAAT tpg|BK006938.2|:957463-958854 7X56=46S 1S1=34S 
 tpg|BK006946.2| 392598 + tpg|BK006946.2| 392696 - INS TTTTGGAACGAATATCTCAATTTTTTAGAGCAGTGGAAGCCATTCAACAAATGGGAGGAGCAACAGCGAATTGACATGCTCAGAGAATTCTACAAGAAAATGCTATGTGTTCCTTTTGATAATCTAGAAAAAATGTGGAATAGATACACTCAATGGGAACAAGAAATAAAT tpg|BK006946.2|:392242-393052 7X6=79S 80S6=7X 
 tpg|BK006946.2| 174563 + tpg|BK006946.2| 175218 - INS TAACACTGTGATTATCAATAAACAAAATGCTTTTCGGATTATTGGGAAATGATAAAATAGTACGAGGTCGGAATGTAGATATTTGTAACATTTCCATTTCTTCTTCCATTTCATCTTCTTCCTCTTCATTGCTTTCATCTCCTCCACCGTTCTCTTGCTTGTTAACACTTGATTCATGAACGTGAAACC tpg|BK006946.2|:174171-175610 7X2=1X144=18S 1S1=165S 
 tpg|BK006946.2| 595110 + tpg|BK006946.2| 594944 - INS GGAATTAATAAAGCCCCAAACCTGTTGCTGGAAAAGACGGTACCACGATCCTAGTTGAAGACCTTTTTTTCAATATTCCTTCTAGATTAAGGGCCTTGAGGTCCCATAATGATGAATACTCTAAAATATTAGATGTTGTCGGGCGATACGCCATTCATTCCAAGGACATTGGCTTTTCTTGTAAAAAGTTCGGAGACTCTAATTATTCTTTATCAGTTAAACCTTCATATACCGTCCAGGATAGGATTAGGAC tpg|BK006946.2|:594424-595630 7X162= 238=7X 
 tpg|BK006938.2| 1486147 + tpg|BK006938.2| 1486426 - INS TAATAAGAGTAGATTTCAATTCCGCCAGAAAAAAAATTTCCTGTGCTAACAGTTCAATGTCTTCGTCGGAATGCTCCAGGTTGACCACCTTAATTGCCACAATTTCTTGCGTAACTCTATCCACTGCTTTATACACATCACCAAAGTTACCTCTGCCAATACATGATTGGATGGAATATAGCTTCGATGGAG tpg|BK006938.2|:1485749-1486824 7X9=1X5=81S 91S5=7X 
 tpg|BK006938.2| 481884 + tpg|BK006938.2| 481312 - INS TCTTCGTCTTGCCTTAGGGATTGTGATAAAGTTGAATATGTCTTAACTTTGAAAGTATGTCGGTTATATGAACTAGGAAGTGTCGCTATACCAGAGGCACAATTTATGGTGGCAGGCTGAATAGTATCAATATCATTTTCCATTTTATCCTTTTCTTCATAACCAGAATCTGCTTTACTTTTGTGAGGATAGTATGTTGCAGAAGAAACAGGCTTTAACGTTAAGTCCTCCGATATTCCATGTAAGCTCTCCTGATAAGTGGACTTAGGCGAAATACATCCC tpg|BK006938.2|:480734-482462 7X4=181S 141=7X 
 tpg|BK006938.2| 460279 + tpg|BK006938.2| 460556 - INS TTTGAACCCATCTAATGTACTGGTATCACCAGATTTCATGTCGTTTTTTAAAGCGGCTGCTTGAGTCTTAGCAATAGCGTCACCATCTGGTGAATCCTTTGAAGGAACCACTGACGAAGGTTTGGACAGTGACGAAGAGGATCTTTCCTGC tpg|BK006938.2|:459963-460872 7X7=68S 71S5=7X 
 tpg|BK006938.2| 419993 + tpg|BK006938.2| 419813 - INS ACCCACCTAGTCGTTTCAATGGGATGATTGCCCTTTAAGCGCCACCTTGTTGTGCCTGTGATGCCACCTAGCAACTCGAAATTCAGTTTTTCTGAAGAATCGATGTGTAAGCGGCACGTCGAAACTTTTAAAGTACCACGAGGCCTATCAAC tpg|BK006938.2|:419495-420311 7X5=71S 71S5=7X 
 tpg|BK006946.2| 442251 + tpg|BK006946.2| 442030 - INS AAGAGAAGCATTTGATATGCTTTTTTTTTTTTGCCGTTTCCACTGCAATCAATGGCGATATAATCGGATGAACAATAAATATTCGTGTTCCTATTCGTCTTCCTATACGTGTTCCTAGCAGCAAACAATAACAGAAGAGAAGCATTTGATTTTCGTAAAAACTTCAGGTGTGGGTGTTTCTTATTAACGGTTAAACTTTACGAATTGAATCCCCTATGTATAATGGTCCATAATACATCTTAAACCACCAAGCCATCTTCGTAATTTTGAACTGGGAAAATTGGGAAAACTGCAGACATTCATAATCATGACAGGATCTTTAAACAGACACTCACTTTTGAACGGGGTAAAAAAAATGAGAATAATATTATGC tpg|BK006946.2|:441270-443011 7X48=1X112= 112S238=7X 
 tpg|BK006938.2| 41384 + tpg|BK006938.2| 40834 - INS CATCTAGTTTGTTTGTAGACACTTGTTATAATGTTCCATTAACTCTGCATTGCCACTATGTGGTGATACACATACAC tpg|BK006938.2|:40666-41552 7X6=20S 58=7X 
 tpg|BK006946.2| 553968 + tpg|BK006946.2| 554115 - INS GGACAAGGCCTCTGCTAAAATATCGATAAAAAAAGAAATAATATGAAAGACAAAACAAACTAACTGGAAAAAATAAAATAAAAAACAAAACTGATCATCATTTAAAAATGTTATTCTCTTGTATCTATTTCTACTAGATAGATGAATCTCTACCCAAGAAATAAACTTTAGCCCAATCCATAGCGACAAGAACTCTGTTTCTAAAGGATAGAC tpg|BK006946.2|:553528-554555 7X5=101S 101S6=7X 
 tpg|BK006938.2| 743948 + tpg|BK006938.2| 743556 - INS CCTTTTGGTCTATCACGAAAAGATAAAACAAGAGCACCGTCGGGTTGATGGCCCCCATTTCCGATGCCAAAGCTGGGCCCAGTACCGTTGGCAATCGTGCTACCGGATGCTGCGCTGTTGTTTTCGTTATTATCATTATTAGATATATTGCTCAAATGTGCTAATCTCTCCGGAGTGAAATAGGAATACTGAATGGAAACGGTTATGTTTCTTGTTTGCTCAGCACCACCATTGAGTGGACCGGAAGCTGCATTTGAATTATTATTATTTTCAGCATTATTTGGTGATGTATTTGTGCCTCTGTTTTGTTCTTGACCACTTTCACTCATAATGAACAAAAGCTGAGGTTACAAG tpg|BK006938.2|:742834-744670 7X7=294S 332=7X 
 tpg|BK006938.2| 1053489 + tpg|BK006938.2| 1054068 - INS GAGGATTTGATCTTTATTTATTGTGGAATCGACCGTAGGTAGATTAGGGAATTTGTGTTTCTCATTATAAAGAGATGTACCGGAAAGTCTCTTGGTTCTGAATTTCTTGCCTAATATTAAACCTTCTAGCAAATCTAATTCCTTTATGCTGTGTGCGATGATGGCACATTTTATAACTTCGTTTGGTGAGCCCTCTCTGTCTCTAAAGCATATCGAATTAATGAGCTGGTTGAGAACTTGAAACTTGTGGCTCCCAGCAATAGAGCTTTCCGTGGGCTCCATTCTCAAAAGC tpg|BK006938.2|:1052891-1054666 7X6=2S 274=7X 
 tpg|BK006938.2| 1071091 + tpg|BK006938.2| 1071478 - INS GAGTAGAAGCAGTGGAAGTGTCCAGAAAGCAGTATGTTCCTAATAATAAAGGTAGTTCTTGGTCTGTGTGATCCCAGCTGGTCAACAAGACCCACGTTGGTCAATTGAAATACTCTTGTGAAGTTGTGCCAGAAAAGGGCCATAGGGTAACATACTCGTTCTATGTGATAATCAACTGTTATAAGCACTATATAGTTACATAGCTGGCCTATACATCTCCTGAATAGTGATGCAGTTTAGAGTTCATCGTGGGCTGCTTCGCTAGCTTCCGCTTTGATCTCTTCCTGTAGCTTGGCGGCGTCTTTATTGTCCAAAGG tpg|BK006938.2|:1070443-1072126 7X142= 159=7X 
 tpg|BK006938.2| 355410 + tpg|BK006938.2| 355506 - INS CATAAATAGGATCTTTTTTTTTTTTATTTTTCATTTTCAATTACAAACTAAGACATAACAATAAGCAGTGCTTTTTCTGTGCATGTTTTCCTCTTTTTATAATGATATTGGCTAAAATAAAATTAACAAAAACAGATGAGTGATATAGATTATATTCATTACAGTTCGTTTTCCTAACTCACATAATAATAGCTTCCTTTGGAACATTATCGGAGATAGACTTATGAGGTAAGACTTTACCACCGTTGATGTAGATTTCGTCCTTAACTTCAACGTCGTCACCCAAGACAGTGACAC tpg|BK006938.2|:354802-356114 7X165= 42=1X236=7X 
 tpg|BK006938.2| 1277995 + tpg|BK006938.2| 1278215 - INS AGGCCCTGAACAGGTACATAGAAGATCTACATTAGAAGGTTTCCCATTCCACCCCTTCGTTAACCCACACGCAAATACCCAGATAAGCATCTTGCACCCCTCACACTTGTATATACGGAGCAAACTACATAATCTCTAAACAGAAAAAAAAAAAAAGAAAGAAAATTAAGAACATTACTTTTTCCGAGCAACAAACGCAAAAATATATGAAGTGGCTGTAGAACAGGCCTTACGGAAGAAAAGAATGATGATGGCATCCCCTTCCCCTGCCCTGGAAGGTGGCCTGTATTTCTGTTCTTTTTTTATTTTTGTTCGCGCAAAGAGCAAGAACATTGGTTGCTTTACTTATTATTTTCAGGGTCGCTTCCGCGGGATGCCATGCACGGATGCCTGCGGAGACAGTGGCGCGG tpg|BK006938.2|:1277161-1279049 7X5=1X142=1X8= 20=1X184=7X 
 tpg|BK006938.2| 491036 + tpg|BK006938.2| 491416 - INS CCTAGGAAGGCTTCTGAGGAATTGTTTAGAATAGATGAAAACTTAGCAGGTATCCTATTGAATTCTTAGCATGTTTATTGTTACGACTAATAGAATTTGCCAGTCAAAATTTACAATATTTGCGTTAATTAACTACAAAACCGGCGGTGCCGAAGGCTTGATAAAGGTAGCACATTTTTATACTGATTCATTACGTTTACGATAGTTGATTGGGTAAAATTTCTTTTTATTTCACTTATGCGAATAACTTACTAACCTTTGTATCATCCTTTTTTTAGCAACCACACATCTTCAACAACCCAAAGGTTAAGAC tpg|BK006938.2|:490396-492056 7X11=17S 294=7X 
 tpg|BK006946.2| 552440 + tpg|BK006946.2| 552760 - INS TGCTAACGCTATTAAAAGATTGTTTGGACTGCCCGTATTTGCTTTATTTTTAAGGACAAATTTAAAAGTCATACAGCAATGGAAGAAAATAAACTTAGTGGAAATAAACCGATTCAACTTGCTACCTGGTCGAACCAGATGGGTTCACCAGAAAACAATGGAAATAATGCAAATAATGGTAGTGATGTACAG tpg|BK006946.2|:552042-553158 7X6=90S 88S8=7X 
 tpg|BK006946.2| 353936 + tpg|BK006946.2| 353549 - INS GGTGCCAAACATTTTTTTTAATCGCTGTTTTGTCTGTTTTTTTCGATTCAGTTATAGGGAAAAAAACGGGAAAGGAAAGAGAAAAAAAAATTAGTGCAGAGCAATAAGAAGCGAAAATCAAAAAAAAGTTTTGGATCTGCAAGACTTGCTGTCACGCAACAATATTATAGCCACCCAGCAAAAATGTCAGACATCGAAGAAGGTACGCCTACTAATAATGGGCAACAGAAGGAGAGAAG tpg|BK006946.2|:353057-354428 7X4=182S 225=7X 
 tpg|BK006938.2| 1268657 + tpg|BK006938.2| 1268740 - INS TGAATATACCGTCCTAGCACTGGGTAAAATGGTGTTTAATCATACACGGTGGCTATTTGGTTTCTATTCCAAATTTGATGTCTACTCTATCGTCGTTACATTCCACCTTGAAAAGGCGTTCCGACTTATTACCAAGGCTACTAGCACTGGATGCAAGGTTAGACTGTACTATAAATAAATTCAAAACTTTGAACTATGAAGCAGGCGACATCCACGCATCCGAACCAGTTGTCGAAGAGGACGAAGACGACGTTGAATATAACGAAGAACTCGATGATGCCGGCCTTATAGAGGAC tpg|BK006938.2|:1268051-1269346 7X170= 2S195=1X80=7X 
 tpg|BK006946.2| 51702 + tpg|BK006946.2| 51793 - INS CATCTCATCTTCATCCAAGTCTTTAGATACAGAAATTCAGAATGTGAAAAATTTGAAGCGATTGTCGATTGGTTCAATGGATTTGGTAATTGACCCTGAGCTAGAGTTCAAAGTGAACAGTAGAAACTCATATTCTTCAGATTCCTCAAAGGAATCCCTTCAAGAATCGCTCCATGAAGAGAAC tpg|BK006946.2|:51320-52175 7X5=146S 161=7X 
 tpg|BK006938.2| 844379 + tpg|BK006938.2| 844400 - INS ATCCAAAAGAGGTTGCGTTACCATTGCTCTTCAAACTTATGTTCGGATCTGTGTTTGGCATTGTTTGCCCAAATGAAGGGTTCGATTGCGAGACTTTGTTGGCATCGTTTTGTGGTGTAATTCCGAATGAAAAACCTTTATTACCAAAAGAAGATTGAAAGTTGCCATTGGTATTTTTA tpg|BK006938.2|:844007-844772 7X7=82S 85S5=7X 
 tpg|BK006938.2| 955559 + tpg|BK006938.2| 955291 - INS GTTTGTATAGTGTAACCCAAAAGG tpg|BK006938.2|:955229-955621 7X4=8S 12=7X 
 tpg|BK006938.2| 1322147 + tpg|BK006938.2| 1322347 - INS TATATACATATAACCATGGTGATGGTATTTTGTTGATAGATAGCGAAATTGCTAGAACTTACCTGTTAAAGAACGACCTCGTTAAGGCAAGAGATTTATTAGATGATTTGGAAAAGACATTGGATAAAAAGGATTCCATTCCATTAAGGATAACAAACAGCTTCTATTCTACAAATTCCCAGTATTTTAAATTTAAAAATGATTTCAATTCTTTCTACTACACAAGTC tpg|BK006938.2|:1321677-1322817 7X12=10S 200=7X 
 tpg|BK006946.2| 624837 + tpg|BK006946.2| 625455 - INS TTTCTTTTTTTTTTTTTTTTTTTTAATTTTTTTTGTGTGGGGAAAGACCGACTACCAGTAATACTTTAAAGATATTATTAAAAGAAATCCCGAAAAAAGAAAGACCATGAGAAAACCGAGTGCGTTTCATGCATGTAACATAATATTTCTTCCCCTCGTTAAGTG tpg|BK006946.2|:624493-625799 7X95=28S 1=160S 
 tpg|BK006938.2| 138785 + tpg|BK006938.2| 139541 - INS CAGTAGAAGAGTGCATCGACATTCATAGATCTCTAATAACATATATTTAAGTGGATATACGCAAAGAAAGGACAAGAAAACTTGTTTCGGTAACAGCATTATTAATTCTGAAGAAATACGCACAAAGAGATGATTTCTGACTACGATGCTCTTTTGCAATTCAACAAAAAACCTGTTTCGCAAGAAATGA tpg|BK006938.2|:138391-139935 7X5=90S 85S9=8X 
 tpg|BK006938.2| 1041663 + tpg|BK006938.2| 1041408 - INS GGGCGCATTCTTGATGGTTACAGAAGTCATGTCTTACAGGGGCGGTTATTCTGCTTCCGACAGACGTAAAATAGAACGTGAGATGTTTCACGGAAATTTAAAGGCTGTCATATCTACCAATGCTCTAGAACTTGGTATTGATATCGGTGGACTAGACGCAGTCTTGATGTGCGGTTTCCCACTATCAATGGCGAATTTTCATCAACAAAGTGGTAGAGCTGGAAGAAGAAATAATGATTCTTTAACCCTCGTGGTTGCAAGTGACT tpg|BK006938.2|:1040862-1042209 7X5=5S 26=1X223=7X 
 tpg|BK006938.2| 610518 + tpg|BK006938.2| 610287 - INS GTCGATGTTGTTCTAACAACAAAACCACGAATCACACCAAAAAGAAGTATGTAAAGGCATGGAAAAAGAAGTAAGCATTGGAATATATGAAATCCTGCTTGTTGATATTCCATTTCTGTGCGAAAAAAGAGCAATAAGCTGGCTTTTAATAATGGGTTGGAGCCATGGATAAGTACGGACATATAGCTCATCAAGAAGGCGATGTTTGTTATTATATTCCAAGGCTGTTCAAATACAACAGTTATTATAG tpg|BK006938.2|:609773-611032 7X7=5S 235=7X 
 tpg|BK006946.2| 133116 + tpg|BK006946.2| 133257 - INS TTTTACTCGCTAGACGGTCAATTGTCACAGATCCAGTCAATTCAAGTCTCAAAGGGTTTGCCCTTGCTAACCCCTCCATTACGCTGGTCCCTGAAGAAAAAATTCTCTTCAGAAAGACCGATTCCGACAAGATCGCATTAATTTCTGGTGGTGGTAGTGGACATGAACCTACACACGCCGGTTTCATTGGTAAGGGTATGTTG tpg|BK006946.2|:132696-133677 7X7=5S 11S180=2X5S 
 tpg|BK006946.2| 106361 + tpg|BK006946.2| 106339 - INS AAGAAAACAGTTGAGAAATTTAATTATTAAAGAAAACAATCTAAAGTCTAATCTCTTTCCCACTGTTGATGAACTGAATCATTATGTCGATTTATATCAAGTGGAATTTCATAAATATTTCCCCTTTATTCATTTATACTCAATTATACCATCCAGTGAAAACTATCCTTTAGTAATATCCATCAGTATGATTGGTGCTCTTTACGGATTTCATTCCACACATGCACTACTATTGTCGAAAATAGCAAGGACGAGAGTTAGAATG tpg|BK006946.2|:105795-106905 12S190=36S 30S4=7X 
 tpg|BK006938.2| 132402 + tpg|BK006938.2| 131715 - INS TGGTAGAGACTCCCCGGCGGAGACAGCCGTCAAGTCCATCCATCCAAAAGTGGAGGAAAAACAAGAAAATAAAGCTATCGAACAAGGAGCGTTGAAGTAAGAAAAACAAACGAAGAACTGAATAAACACAGCCTGCTTCAAATTATGGAAGGAGCTGTTACAC tpg|BK006938.2|:131375-132742 7X264= 143=7X 
 tpg|BK006938.2| 318014 + tpg|BK006938.2| 317392 - INS CAATAGAAGCTCTTCTTGCAAAAAATTCAGAATCAGCTTGGAGTTCCTATTGGAATCGTATATGGAGACTAACTTGCTGTACAAGTACAATAGAAGCTCTTCTCCCTTTGTCGAATCACTTTGGTACACGTCGTTACAGTAACTTGTCGCCGCTTTGTAATCATCTATCTCATCAAGTAATATAT tpg|BK006938.2|:317008-318398 7X7=151S 65S97=7X 
 tpg|BK006938.2| 738558 + tpg|BK006938.2| 738666 - INS AAACGCTCCTTTTAATAAGAATATCATTTTCATCTTCTAAACAACCGACAAGGCATCGGATAAGTAGACCTGGTTCAGGGGTTACTAAATCTTTGGCAGCAGGCAATAAGACCTTGAAAGCTTCTTCTTTTCTTTTTTTCCTGTCTAGATGAGAATCGTTGGTTTCAGT tpg|BK006938.2|:738206-739018 7X8=76S 77S8=7X 
 tpg|BK006938.2| 1399011 + tpg|BK006938.2| 1398335 - INS GTCCCTGGTTCTCAGCCATGCTGGTGTTAAGTGTTGAATTTTCCACCGTCTCTTCTAGAGGAATAGTTGTTTGAGTAGATTCCTGTATTCTTCGATCAAAACGCAACTTCAGAGCATCAAGTTGCTGTTTTATATTTTTAACTTGTGCTTCCCTACCACTCACGTCTTCGTTTTCATCCCTTTTCATTACGATTATGCTTCTGTCCAAATCAACTATTGTTTCCTCAACAT tpg|BK006938.2|:1397859-1399487 7X8=68S 116=7X 
 tpg|BK006938.2| 744658 + tpg|BK006938.2| 745230 - INS GGTTAGGGTTGTTATCACCATAGGCGATCGAAAATTCTGTATTATTGGAGTTGAATGTAGACGACTTAGAGGTATTAAATGTCCCGTATGTAGCGCAGTCAATTAACTGTGATGTAGAAGCTGTACTATCAAAAGTAGCAGTGGCTTCGCTGGTAACTATAGTGGTGTCGTAGCTAATTTCAGTAAACACACTCTCAACCACGCTAGCCAAAGCATCCTTGTTTACTTGTTTAAAGGATGAGCCAGTGGTATCCTTCTTTTTAGTGGAACAGTATGGG tpg|BK006938.2|:744088-745800 7X6=150S 261=7X 
 tpg|BK006938.2| 704925 + tpg|BK006938.2| 704931 - INS TACTAGATTAAGGTCATACATATAAGTTAGTTCTTGAGAGTATTAAGGTCAAAGCGGAAGTTGTCTCTTCGGATGAACGTGAATCCAGTCTAAGAAACCTTTTGAACTTCGGACATTCTATTGGTCATGCTTATGAAGCTATACTAACCCCACAAGCATTACATGGTGAATGTGTGTCCATTGGTATGGTTAAAGAGGCGGAATTATCCCGTTATTTCGGTATTCTCTCCCCTACCCAAGTTGCACGTCTATCCAAGATTTTGGTTGCCTACGGGTTGCCTGTTTCGCCTGATGAGAAA tpg|BK006938.2|:704313-705543 7X95= 281=7X 
 tpg|BK006938.2| 634224 + tpg|BK006938.2| 633817 - INS AAAAGAAGGTTTAAGAACATTATGTTTGGCTAAAAGAGAGCTCACGTGGTCCGAGTATGAACGTTGGGTTAAGACTTATGATGTGGCCGCTGCATCCGTTACTAATAGGGAGGAAGAGTTGGACAAAGTTACTGACGTTATTGAACGTGAGCTTATTTTGCTTGGTGGTACGGCCATTGAGGAT tpg|BK006938.2|:633435-634606 7X6=11S 92=7X 
 tpg|BK006938.2| 968037 + tpg|BK006938.2| 968051 - INS CCTGCTACATGCCAAGTTCTTTTGCTGTCCAGGTTGTTTACCCAAAACGCGGTAGAGATTTCTTGCTTGCACGAAATCTACATCACCTGGGGATGTTGCCCAATGATAAGGGATAGCTGGCCCATTCCATACCTCTTGGTGTTGTTGAATGGGTCTGTCCTGTTGGATATACGTGTACGATTTATCGTTGGCCAAATATGTAGGTTCTGAGCCGAAGTTGCCGTTAACATTCATCGGTCCATCTCTGATAGCGGGATTGAAAAATTTAGATGCATATGGAC tpg|BK006938.2|:967461-968627 13S82=1X99= 264=7X 
 tpg|BK006938.2| 691821 + tpg|BK006938.2| 691807 - INS GCTAGAGATAGCATACATTGGACCAGCTAAATGGTATGTCCCCTCGCAGAACTTACATTTAGTATCAACCGGAGGCCCTTGCGCAACCGAGTATTTGGTGAATGTTTTGTTGTTCCTACCTTCGCGTTGAGAAATTCTGCCCAGAGGTTGATTGTGGTAAGAGCCGCAACGGGAACAATGGTAAGTAGTC tpg|BK006938.2|:691413-692215 17S85= 23=79S 
 tpg|BK006946.2| 805961 + tpg|BK006946.2| 806197 - INS AGGTACGCAGATTTCAAAGTCTCTTTATCAGCGGTTGTAGTGGTAAGCTCAGATCCTCGTATAATATCTTCGATAGGAGCATCGATCTGAGTTTCAATTTGACTTTCTTCGTCAAGATCACTCATCAAAACCCCACGTAATGTTTGTT tpg|BK006946.2|:805651-806507 7X5=153S 74=7X 
 tpg|BK006946.2| 609737 + tpg|BK006946.2| 609657 - INS TTTTCTACACTTTCCACCCTCAACCTAACAGAGCCCGCTGGCACAAATAATCGATAGTAGGACAACAGAGCTACTCCTTCTTATGCCCCGCCCCTTTGAGCTTGTTGTATTGCTCTTGATAGTTGTGTTTTTCACTTTCATCAGCATCGGTAGTCTTGCCGTCCTTGTCTTGACTAGCCATTTTCTTAAAAGCGTCACTCACTACC tpg|BK006946.2|:609231-610163 7X75=28S 1S1=226S 
 tpg|BK006938.2| 1102339 + tpg|BK006938.2| 1101644 - INS TTATGTAATACATATAATGATGGGTGACATTTTTTGTGTCATTTAGATTAAAAGAAATTTTAAGAAAAATTGACGTATTTAATTTTGATCCGCAGTAAACGCTATAAATTCTTTTTAATATAAATGACAGCTTTTTATACATATAGACCCTTTGAAGAATATTCCAAACTAGAAAGGTTGATCAGAAATGAGTTATAGTGTCAACACGTTTACAGATTACGTT tpg|BK006938.2|:1101184-1102799 12S163= 112=7X 
 tpg|BK006938.2| 421689 + tpg|BK006938.2| 421039 - INS CTTCAGCCATTGAATCATTTGGGCTACATTCAAATCTTTGCACATGTCCAAAGGCTGCTGATGAGCTTTATTCTTGACACAATCATTGATAGACTTCTGGCTAAGAAGGAAACTGATCACATCCGACCGAGATTGAGCAGCAGCCAAGTGC tpg|BK006938.2|:420723-422005 12S14= 4S129=7X 
 tpg|BK006938.2| 128078 + tpg|BK006938.2| 128178 - INS GGGTACCAATGTTTTAATGGCGGATGGGTCTATTGAATGTATTGAAAACATTGAGGTTGGTAATAAGGTCATGGGTAAAGATGGCAGACCTCGTGAGGTAATTAAATTGCCCAGAGGAAGAGAAACTATGTACAGCGTCGTGCAGAAAAGTCAGCACAGAGCCCACAAAA tpg|BK006938.2|:127724-128532 7X4=38S 36S92=7X 
 tpg|BK006938.2| 1234667 + tpg|BK006938.2| 1234071 - INS GACATTTTTTTTCTGCGTTTATTAATACTACATAAAATCTGATATAAAACATATTTAACTGATCAACCCTCTCAACTTGATACTCAAAACAAGTTGACGCGACTTCTGTAAAGTTTATTTACAAGATAACAAAGAAACTCCCTTAAGCATGGCACCTG tpg|BK006938.2|:1233741-1234997 7X4=180S 79=7X 
 tpg|BK006938.2| 1431016 + tpg|BK006938.2| 1430946 - INS CCCAGCAGGATTTTTCTGACTTGATGAAGTCTTGGAAAAATGAACGGTGTTCGCCAGAACTCTTACCATATCCTCATCAGTTGATGAAAAGATTATTGAATCGAATATCCATGC tpg|BK006938.2|:1430704-1431258 7X81=15S 4S1=26S 
 tpg|BK006938.2| 1520093 + tpg|BK006938.2| 1519884 - INS TCTACAGTGTCTGCTGCATATTTCTTGATAGAATTTAGGATGTTTTTTGTACCTTCTAACGCGGGAATCAATAAGTCTTTTTCATATTCGGTAGTATCATAATGAAAAGGAGAGGCCGTGTGTAGAACATACCTAATCTCACGTCCACGTTTCTGCAGAACCTTATCG tpg|BK006938.2|:1519534-1520443 7X110=16S 38S4=7X 
 tpg|BK006938.2| 1113075 + tpg|BK006938.2| 1112664 - INS TATGCCCATTCTTCTTTTATGGTCAAGTTTTCGATCATTAGTTGCGATAATTTCTTTACCTCTGGTTCAGCTTTTTGCCCATCTTCATTCGTTTTATGGCCCTCTGGGTTCAAAATTGCCGGAAGCGACTTCAACGGTAGGATTTTTTCGTTTATGTATGCAGCGGAAGCTATCTTGATCGAATTTTGAAGTTGTCTCTCTAGATGACTTTGAGGTTCTACACTTAAGAGCTGTCTTGTTAGTGTATTATACAAGTTAAAAGAATTGAGTAATTTATGTC tpg|BK006938.2|:1112090-1113649 7X4=149S 263=7X 
 tpg|BK006938.2| 1292103 + tpg|BK006938.2| 1292274 - INS CAGTAGCTGAGTGCCAATTGCCCACCAAAAGAACCCAAGATAACTTGGATGTCTTGACCAGGAGTAAACGCCAGTTTTCACTAAAACATGATCGGACTCCTTCTTGGTCTTCACAATATGAGAAAAGGAATGTCCCGCAGTATGCATAGCAATAGTTCTGGTATATTGTCCCAGAATAACTAGAAGACATCCAAGTACTGTACAAAGCTTGGTAGCTAGAGAG tpg|BK006938.2|:1291643-1292734 7X207=2S 7S1=46S 
 tpg|BK006938.2| 1017409 + tpg|BK006938.2| 1017559 - INS ATGATTGTACC tpg|BK006938.2|:1017373-1017595 7X5= 3S3=7X 
 tpg|BK006938.2| 805046 + tpg|BK006938.2| 805647 - INS TTACTCTTCCAAATTTTTAATATTTAGCTGGGGTTGGGTAACAAGTGAGCAAGGGAAAAAGTGAACATTTTAAGAAGAACAATAAAATAGCAAGAGATGGAATGGTAATGCTTGGCTCTCGAGAAGAGTAGCATAAAACGAGACTTGTTTAAAACAGGATATGACATACTTCAATTCAGCTTTCCCTATCAGCCGCTCGAGCAGTTATATAGGTGTGTTGCCGGAGTAATTTGGCGGAGGCCAACAGTGGCTAGGCGGCAACGCCTGGAACACGCGCGTAAAAGTTCTGGAAGGTTCGCGAATTGAGAACTGCTCAGGGG tpg|BK006938.2|:804392-806301 7X1=2I205=32S 1=205S 
 tpg|BK006938.2| 1419500 + tpg|BK006938.2| 1419929 - INS GTCAGTGACCACAGTGGATACTATTATCTTTGATCTCTTCGAGATCCGTCTCTTTTTAGGACGAGAGCTCGAGTCAGATCCAGGAACAAGACGTGTCTGTTCGCTTGGTAATGTGTGAGTCATCATGCTGCTAATGCGCGTTCAAATAATGTCCCGTATGCTGATATGTAAATGTTTATGTAGCCACTTGCTGGCAAAATGTGGAGCACGAAAAAATATAAACGTTTAGATACACTTCTTTCTTTATATACTAAAATCCCTTTACTTTTCCTCTACGCGCGAAGCTTATCGCTATCGTCAATGC tpg|BK006938.2|:1418878-1420551 7X200= 152=7X 
 tpg|BK006938.2| 332696 + tpg|BK006938.2| 333317 - INS TATGCGTTCCTTTCCTTTATATCCGTCAGGATTAACTTCAAGGACTTCACACAGTTTTTCTATCTTACTAATATTCTTTTTCGTCACCGTGTTTATAGTTCTGATGGGAATATACCTGCGAATCCCAGATATTCGAGCAACAGTAGTTGCAAACACTTTTGTCCTCAACATGTCGAGATTCATTATCTGATTTATTCTTTTATCCTGCTATAAAGAAACCATAGAAGAATAGAAGCAAAGGGGTAGTACGTGGCACCTCCTAAAGGTAATATTGTACTATTC tpg|BK006938.2|:332118-333895 7X256=8S 1=163S 
 tpg|BK006938.2| 1381663 + tpg|BK006938.2| 1381464 - INS CTTCTTCTCTTCCTTTGATACTTTTAAATTCGGCAATTCTGGTTTTGGAAGCTCTTTTACCCTTGGTTTGTCATCCGAAGAATCTTTCTTATGAAGTTCTTCTACAGTTTCCAGTTCAGAAGTTAAATCAGCAGAAGTTGCTTTCCCATCTGACTTAGAT tpg|BK006938.2|:1381130-1381997 7X6=14S 140=7X 
 tpg|BK006946.2| 571945 + tpg|BK006946.2| 572575 - INS GCTCTTCTGACAATGATGATGAGTATAGTACTACAGTAACGTCCTTCATTCATTACCTTTACTAGCAGTGATAAAAAGTTTTGAAAAAAAATGTGCTCCAGGGGAGGTTCGAACTCTCGACCTTCAGATTATGAGACTGACGCTCTTCCTACTGAGCTACTGAAGCTGTCTGTTATGGAG tpg|BK006946.2|:571571-572949 15S82= 70=27S 
 tpg|BK006938.2| 1448695 + tpg|BK006938.2| 1448991 - INS CTTATATGGGAGGATTGATATCAAAGCTGATTTATACTGACCGATTGCAAAGTGTCCCAAGGTTAATTTCTAAAGAGGATATTGGGATGGATAGCGACAAATTCACTGCCCCTATAATAGGTTACAAGATGGAAAAATGGCTTTTGAAGTTAAAAGATGAAGTTTTAAATATTTTTGAAAATTTATTAATGATCTATGGAGACGATGCGACCATAGTAAATGGAGAAATGCTCATCCACTCCTCTAAATTCTTATCCAGGGAGCAAGCGTTAATGATAGAAAGGTACGTGGGACAAGAC tpg|BK006938.2|:1448083-1449603 13S56=1X217= 14S5=7X 
 tpg|BK006946.2| 565284 + tpg|BK006946.2| 565107 - INS GCTCATATATACAGGAGATGGATGGGTCAAGTTGACTTACAAATCCGAACTTTCCAAATCTCGTGCTTTACAAGAAAATGGGATTATAATGAATGGAACATTAATTGGCTGTGTTTCGTATAGTCCGGCTGCTCTCAAACAATTAGCTTCCTTGAAGAAATCGGAGGAAATTATAAACAATAAAACAAGTTCACAAACTAGTTTAAGCTCAAAAGACCTCAGCAATTATAGAAAAACAGAAGGAATTTTTGAGAAAGCTAAGGCAAAAGCAGTTACTTCAAAAGTGCGCAATGCAGAATTCAAGGTTTCCAAGAATTCTACTTCCTTCAAAAATCCACGCAGGCTTGAAATAAAGGA tpg|BK006946.2|:564379-566012 7X141=1X293= 179=7X 
 tpg|BK006938.2| 1215172 + tpg|BK006938.2| 1215577 - INS CTATCCTCATTTTTCCCC tpg|BK006938.2|:1215122-1215627 7X9= 5S4=7X 
 tpg|BK006938.2| 864502 + tpg|BK006938.2| 864714 - INS TAGTAACAATATCTCTTTTTTTTTTTCAGTGAGCTTTTATTTTTTTTTCATTGCTCTTCTTTTGGCCTCTTTTGTTTTTTTCTTGATTTCCTCCAGTTTCATCTGTTTTTTCTTTGGATCAGATACAAAATCTGGTTTGAACGCGTCATAGTGACAGTCCAATTTCAACCTTTCACAGTTGAAACAGTGCGGTCTTTCCTCGGTACACTTCTTTTTCCTTAATCTACAAATCCAGCAACCAGTACGGGAC tpg|BK006938.2|:863988-865228 7X125= 11S3=7X 
 tpg|BK006938.2| 33676 + tpg|BK006938.2| 33996 - INS CAATATTGATGTATTGATGATTATGTGGCATAAACGAATTATATCTCCGGTATTCAATATGTAAAGTTCCGTTTCTATTTACCACTATTTAACGGAATTTTTGCTCCTTTGCCCTTCATGTCTTATGATAGGTTTTTTAGAAAGAAGCAGGGTCAACCTCTCGCTCTGACAAGGCAATACGCCGGTAGAGGATGAGGATGAAGAGGAGGATACGTTTTGTAAATCTCTTTCCATGACGTGCATCATTTTCTCAAACTTCTTGAACAAAAGCTCTGCTCTAACC tpg|BK006938.2|:33096-34576 7X10=1X166= 142=7X 
 tpg|BK006938.2| 263765 + tpg|BK006938.2| 263387 - INS AAAACCATTCAATGCTACTGATCTGATAGGTGATGTAATCTTACCATTAGACCAGGAAATGATTAGGCCATTATTGGCCACTTCGCTTTCGTTGGCTGCAGGGTCCAATAGCATATTGTTGCCTACAACGGCCAATATAAACACTAAAGGCGGATTAATGTCAAGCTTAACCATGTCGTAATCATGAAACGTAGGAAGTTCTTCCACCTCTAAGTCGTCAAAAGCTGAAATAAGTTTCGGTAGGTATGTGGAGTTCAACGC tpg|BK006938.2|:262851-264301 7X4=212S 131=7X 
 tpg|BK006938.2| 270215 + tpg|BK006938.2| 270226 - INS GTAGTATTGATCGTAGGTAATATTTCATTCGATGATTTATAGTCTAGAATTAGAGAATTCATGAATCTTAATGATTTCTGTAAACCTTTCAAAGTGTGAGGAATATTCGAACCACCAACAAATGCGTCATTTACCTGTCTAC tpg|BK006938.2|:269917-270524 7X7=64S 68S3=7X 
 tpg|BK006938.2| 783769 + tpg|BK006938.2| 783785 - INS TCTGTACTTAGGTAGGAATCAATCAAATCAACAGATGTGACATTATTTAAAAGTTCTTGGGGTGTGAGGAAAAGATAACTCAATATTGTCTCCACAGTTTTATCGATAATAAGAAACTTCAAGTTATTTTTCGTCTCAATCTGATTCAAAACCCCTATCAAAT tpg|BK006938.2|:783429-784125 21S67= 23=66S 
 tpg|BK006946.2| 278917 + tpg|BK006946.2| 279168 - INS GTGTTCGTCATGCACACACCACTTGGCCATGATTCATCAGTATTGTCGGATATATCCAATGCGAACACCACATCCAAGTCACGTTCCTTCTTGATTAGTGGAACCAACGGCAAATTTTGGCCGTCCTCACCACCATCAACTAAAAACAAATCATCGGCATCAACAAT tpg|BK006946.2|:278569-279516 7X4=79S 79S5=7X 
 tpg|BK006938.2| 47352 + tpg|BK006938.2| 47626 - INS TGATAAACCGTAAGGTTTTTTGGAATTAT tpg|BK006938.2|:47280-47698 7X4=10S 15=7X 
 tpg|BK006938.2| 1204524 + tpg|BK006938.2| 1204632 - INS GTTATTTATTGTGCCCTGAGTTTCGGTATCATCATCATCATCCATTAAAAGCTCCAATTCAGCCTTTGATTTGGCATTCTTTTCGATCTCCTCTTCATCGTTAGTATGC tpg|BK006938.2|:1204292-1204864 7X6=48S 51S4=7X 
 tpg|BK006938.2| 284000 + tpg|BK006938.2| 283523 - INS CCACAAACTCAAGAAGCTAAGGCAATGAAGAATCTGACTTTCTCACCACAATTAAAAAGCAAAAAGAAGAAGATGAGTTGACCAAACTAAGGGCGGAAAATGAGAAACTCACACAGGAAAATAAACAACTGAAATTTTTGAATATGGAAAATGAAACTACTGTCGATGAC tpg|BK006938.2|:283169-284354 15S151= 28=1X120=7X 
 tpg|BK006938.2| 425857 + tpg|BK006938.2| 425202 - INS TGTTTATGTACTATTTTTGGTTGGAAAGAATTAAGAAAATGCGCAGCGTTGCATGGATTGGGTTTCGAAGCTAGTGGGCTCATTTGGGATAAACCAAACGGATATTCTAATGGATTGAAGGAATTTGTTTATGATTTGCTTAATAAAGAATGTACCATAGGTACGTTCCCTGAGTACAGTGTTGCTTTTGAAACATTCGGATTTCTACAACAAGAATTACATGACAGGATGTCCATTGAACCTCAATTACC tpg|BK006938.2|:424686-426373 7X4=7S 126=7X 
 tpg|BK006938.2| 1069498 + tpg|BK006938.2| 1068786 - INS CTTCCGAATTTGCGTCGCTATCAACAGGAGCTGCTGCGCCTAAAACTCCATTAGAAACTGTGCTATTTTTCCTCTGTTCATAAAAATCCGTTTTTATCAGAGATTCTGAAATTTTACTCAACTCGTGATTTAATTTAATCAACTGCTCTGCAGATATGCCAGAAAATCCGTTATTAATGGAATAATTTGAATCGGCGCTAGTCGTTACCTTATTCTCCTCAAGATTTTTGATATACTTGGAGA tpg|BK006938.2|:1068286-1069998 14S17= 122=7X 
 tpg|BK006946.2| 532162 + tpg|BK006946.2| 532672 - INS CCACCATTCTCACTAACTTATGTAAGGACAGAAGAGACTGATGGAAAACACGGCAAAAGGAGGTCGCAGGTTGTTGAGACGCATAAAGTCACTGATATATATTCTCATGAATACAAGGTAATTACAAGCTTGCAAGGTACCTACGAGGCGATTGAAATTACAGATGCTTATTGTTTTGCCA tpg|BK006946.2|:531786-533048 7X4=86S 86S5=7X 
 tpg|BK006938.2| 1475524 + tpg|BK006938.2| 1476153 - INS AGTGTAGCAGTGGGATTCAACCCCTTTTCCATACATTCAATGAAGTACGCTGTTAGTTCGTCCAACTTTGCTGCATCAACCTGCAATGAGGAGCAG tpg|BK006938.2|:1475318-1476359 21S27=7S 43S5=7X 
 tpg|BK006938.2| 500550 + tpg|BK006938.2| 500563 - INS TTGCTAGATTTGTTGACATTTTTGGATTTTTCTTATCTCGTCTTCGTCAATATGCTTGCTTTAGGATTTATAATCTTCAAGGATATTATCTTTTCCCCCTTGCTTTGACTTTTCAACGTTCGTACAGAACACCAGGTGTGTGGTTATACGTATAAC tpg|BK006938.2|:500224-500889 7X29=49S 3S1=246S 
 tpg|BK006938.2| 494153 + tpg|BK006938.2| 494263 - INS CCTTAGAGAATATAACATCGATGATTCATTAGTTTAAAAAGTAAATAATGGTACATAGCTTGAAATCTAATTTTTCTTTATCATGTTTATACAGGCGGAGGTGGGGCATTGGCCATGTATATTTTATTCGATGAGGCCTGGAATTGCCCCAACAGGGTTGTATAATGA tpg|BK006938.2|:493803-494613 8X50=33S 5S1=15S 
 tpg|BK006938.2| 656709 + tpg|BK006938.2| 656701 - INS CATCCCAAGTCTTGATGGGACCTAGTAG tpg|BK006938.2|:656631-656779 7X2=12S 12S2=7X 
 tpg|BK006946.2| 902942 + tpg|BK006946.2| 903643 - INS GTACAGCTATTGGCGCAAGAAGCCAAGGGGCAAAGACTTATCTAGAGAGAACTTTAGACACGTTTATAAAAATTGACGGGAACCCGGATGAACTAATCAAAGCTGGCGTCGAGGCTATCAGCCAGTCTCTAAGGGACGAATCCTTGACTGTAGACAATCTTTCAATCGCCATCGTGGGTAAGGAT tpg|BK006946.2|:902558-904027 7X6=86S 89S4=7X 
 tpg|BK006938.2| 600838 + tpg|BK006938.2| 600498 - INS AAGCTCCAACGTCATGCGGCAGCGTCAGATGTGTTAAGAGACAGGTGTATTTTTGATTGAAAATGATTTTTTGTCCACTAATTTCTAAAAATAAGACAAAAAGCCTTTAAGCAGTTTTTCATCCATTTTACTACGGTAAAATGAATTAGTACGGTATGGCTCCCAGTCGCATTATTTTTAGATTGGCCGTAGGGGCTGGGGTAGAACTAGAGTAAGGAACATTGCTCTGC tpg|BK006938.2|:600024-601312 7X4=217S 16S186=7X 
 tpg|BK006938.2| 446035 + tpg|BK006938.2| 446022 - INS TCCTTATTGGTTTGAGTT tpg|BK006938.2|:445972-446085 7X5=4S 7S2=7X 
 tpg|BK006938.2| 627399 + tpg|BK006938.2| 628088 - INS GTTCTGACAG tpg|BK006938.2|:627365-628122 7X5= 5=7X 
 tpg|BK006938.2| 1114909 + tpg|BK006938.2| 1115286 - INS TTGATCCCTTCGCAAGAGCATATGACAATTTTGGAATTATCGATGAACTTGACTAATTTTGTGGAAGTTCTCAATAATAGGTCATTATCTAGTTTAGTCACTTTCAATTTATTACCTACGGGCTGTAAATGAAAAACTTTAGTGGTAGAGGGCCTCCCTACGACTAAAACTTGTCCATCAGGTGATAAAGAACAAGTTGAGATATTCTGGTCATCTTTTAAAGTTAACTTGCAAACTAGCTTATAATTCTGTTCTGTACTAGAATCGGTTCCCATTGTC tpg|BK006938.2|:1114337-1115858 7X7=10S 140=7X 
 tpg|BK006946.2| 886134 + tpg|BK006946.2| 885622 - INS CTGCTCTTCACCGCTTTTTCTTTCATTAATGCACAAACAGGGGTCTCTGACTCAACACCAACTAGCGCTGTTTTCCGTTTGTTGCTCGTAACTTTTTTGCCAATCTTTCTTAACTCAATAGTGCTTTTTCTATTATTTTGGGTTTCACTTTTTGTGGTTCCTGGATTGTCATATTGTTGTAAAGACGCAGGTGCCGTGATTGCGTTTATTGCACACACTTTCTCGGTTTTGGGCTATCTTTTAGATTTCGAACTGATGTGGTTCTTACAAGGTTGGAACTTTACCCGTACATTGATACTGCTTATTACGTGCATCAATATGCATCTGATTCTTTTCAAGGTCTTTACGACGATATTCTTGACAAGGGAGTATAAAAACAATAAGGCACATTTGGCATGGTGGAATGG tpg|BK006946.2|:884794-886962 7X5=160S 29=1X174=7X 
 tpg|BK006946.2| 409584 + tpg|BK006946.2| 409956 - INS CAATGGCAGCAATGGCAGTTAACGATAATAACGGATCAATTTCAATTCCAACTACAACAAAACCCTTCTCCAAATTTGAATCTCAATATTAACCCGGCACAACCTCTGCATCTACCTCCTGGTTGGAAAATAAACACTATGCCGCAACCACGTCCTACGACAGCACCTAACCATCCCCCTGCGCCGGTGCCTTCTTCGAACCCTGTGGCCTCGAACTTGGTTCCTGCCCCATCATCAGA tpg|BK006946.2|:409092-410448 7X169= 6S219=7X 
 tpg|BK006946.2| 653851 + tpg|BK006946.2| 654046 - INS ATGATAATCAAAAGAAAAAAACAATCTACCTACATATATATGCACTCAACATACATAAATACACACGCATTATTGTTTCTATAAACTTCCAACAGACAATATTCCCATACAAACATCAACTAACTGATTTCCTCTTCATACGCGTTCGCTTCACGTGATGTTCCTTTTCCATTGAAAGG tpg|BK006946.2|:653479-654418 7X4=85S 86S4=7X 
 tpg|BK006946.2| 415306 + tpg|BK006946.2| 415873 - INS ACAGATTATGACATGGCATTTGGATTAACGTAGTCGTGCCGAACGAACTAGATTCTATACAATTCAATGACTTTTCCAGCGATGAAATAAAGCATCTGTTATATTTAAAGAAGATTATCGAATCCAAACCAAAGGAAGAACTGTTAAAATTTTTAAACATAGAAAATCCCGAAAACCAATCCGAATAGAAACGGCGTACATACATAAAGAATAAATCAGGAACGTGAACACCTTCCTTACATATATACACACATACATAGGCATATGTATCGCATCTTAAAGTGAGAGATCTACCTATTTTCCTTTTTTTTCCATTTACAACATAGCAATTGATGTTTTTTTCCCTTCTAAGTCATCTCGATGTCATCATCTTCATCGTCTTTGTAGTCAACTTCTTTCCTGACCCTCAATTTCTTCATCACAATATTTT tpg|BK006946.2|:414432-416747 7X320= 12S405=7X 
 tpg|BK006946.2| 607251 + tpg|BK006946.2| 606572 - INS GGGCGTATGTTATAAACCTAAAACAAGATAACTATAAAGTTATGAACAAATTGAATATATTACTTAAGTTGGTTGCGCAGCCAAGCGCGCGCCCAAGCACAAACAATGCCCAAAATAAGCTTGCTATCGAATTGCTAAATTCGATATCAGCCGTTAGTAGTGCTTACTTGCAGAAAATGCAGAATAATGGCTCTGGTAGACAGCATACTGCTGATTTATGTACAGGAGATTCCAACACCCATTCTGGTATCAACCAGCATCGGACTACGAATGGAACCATAGATGTGAATACGAATACTGCAC tpg|BK006946.2|:605952-607871 7X5=152S 285=7X 
 tpg|BK006946.2| 755230 + tpg|BK006946.2| 754770 - INS TCCAGAGCGGTATGGGGGTATATAGTTTATGTTCTCTGTAGAACCATGGGATAAATTCACCGACGGCTTCAGCCCTTTATATCTTTATTACAGGCAATTGGAAGTATTGCAGTTTACAGCGTCATCTACAATACAATTAGATGATGCTGTAGTAGCACCATAGGCAGTAGGTGAACGCTTTTTTCTACCATGCTCAGTGTTTCCATGGCTGTCAAAGGCTTCTTGAGACGAAGATGGTGAACCACCTGCTATGATAGAAAATCTTCTGCGAATATCCTCATTAACATCTCCAGAAACAAATTCTGGTTGAACAGTTGCAGAATGAATACCGTGTTGATGGAATATTTTTCTTATCAGCTTGGCGGAGCTCATGAATTTATCAGGTGCACAGTCTATTTG tpg|BK006946.2|:753958-756042 7X6=5S 5S382=7X 
 tpg|BK006946.2| 669542 + tpg|BK006946.2| 670012 - INS TTTATAGTCGATAAAAGGTTATGAACTATATCTTTTGTTTTGCTGTTTCGAATGAATACTTGGGGCTGCTATTGGAATATTCAGTACAGGAGCGGTTCGTCTGATAGCATTTTTGAAAGCTTCATTTATGGAGATTGACACGGCATCGGTAGGGTCGCTCGGATAGAGAAAGCTTGCATTTAGATTAGAGCAAGTGTTCGATATCACGGAGAAGCTATTATCTGTACATCCTTGTTCGTATTCTTCATCCAGCAAGTAATTAAGGTCGTCATCATCATAATTA tpg|BK006946.2|:668962-670592 7X8=178S 142=7X 
 tpg|BK006946.2| 810921 + tpg|BK006946.2| 811572 - INS CCTCTTTCTTTTCTATCTCTATTGCGCCTTCCAATTGTGGTTGTAATGGTATCTGCTGCTGCGGCTGAGAATCTTTAAGGGTTTTTACGCTTATTTTTTGGGAACCATGACGGCTGTGATGGTGACGGTGAGGACGAGGGCGATTGCGCAACACAATGGGTTCAACCGGCTCCCTTCCACTTTTGTTACCAAGCTTTTTGCTTTTCCTCACGCGAACGTGCACGGCATCGTTATTTGGTATTGATGGTGACGATGATGGTGACGACGAGGGTGATGATGATGCATCATGCTTGTGGTGTGGCTTTCTTC tpg|BK006946.2|:810289-812204 7X289= 45S4=153S 
 tpg|BK006946.2| 431548 + tpg|BK006946.2| 431090 - INS GTGTAATTGTATTTATAATAGTGAGTTTCGGAACTTAAAAATCCGTTTCCCCGTCAAGAGAAGCAAAGATCAGTTCATATAGTGATTTCCCTTAAAAAGTTACCACAGCTTCTGAATTAACTGTAATCCTTATCTACTAGTATCAACCAACCCTTGTGTTTTTTTTTTTTTT tpg|BK006946.2|:430732-431906 7X86= 175S5=7X 
 tpg|BK006946.2| 319532 + tpg|BK006946.2| 319080 - INS TACTATATTCTACACTCTCACCTGGTGCCAACATTGATGCTTGCATCTTGTGGAGAGATAATAGACCTGAATTTGAGAGACAGGTAAAGTTATCCATTTTGAAATCATTAGGATTCTGAAAGCAGGTAGCAGGTTAATGATCATTTGGTCTTCCTTTTAACTGTTCTCTATATACATAAATAAGCATATCTACCA tpg|BK006946.2|:318676-319936 7X3=177S 10S173=7X 
 tpg|BK006946.2| 575239 + tpg|BK006946.2| 575987 - INS TGGATTGGCTCTTGTTCAATTGGGATACGTTTCGACTGACATTTTTTGGTAAGCTTTATGATAATTTTATGACAATTTCAGAAAAACTTGCTATAGATTATAATCACCCTAAAATCTTGAGAAATTTATGGTGCAATGGGAAGTACATGGGCATTGATTTAAAGAATGCTAATAATTTAAACCTTGATACCGATGATGAAGCAACTAGTAACATTAATGA tpg|BK006946.2|:574785-576441 7X10=100S 102S8=7X 
 tpg|BK006946.2| 271743 + tpg|BK006946.2| 271448 - INS TTATTGATGCTACATAGGCTTTGAAACTGCCGCTTGAATTGGATTTACTTTCTCAGTGATTCTATATGTATTGTACGAAAGTTGAGTAGCACAAGAGTAACTGTTCAAGATATGCCTTGTTTCAAAGGATGTACATTCAAAGATCATCCCAGGTCCTCGAGATATTTATTCGTTCTATATTTTGGATTTTCTTTATTGGGTTTGTTTTGTTT tpg|BK006946.2|:271010-272181 103S10=119S 5S194=7X 
 tpg|BK006946.2| 512365 + tpg|BK006946.2| 512455 - INS TTCTCTCCTCTGTCTTTCTTTGCCGAGCTCCATCGTGCTAGCGCATCGGACAGGAAGCAGTGAAATACAAGAAAAGTATACGAGCAGTATTCCTGCTCAAGAACCCAGTTTTCAGTTATAGTTTCCACTCCTTTCAATAGATGGGAAACTATATATCC tpg|BK006946.2|:512035-512785 7X4=75S 74S5=7X 
 tpg|BK006946.2| 215270 + tpg|BK006946.2| 215499 - INS ATATGTATGGTATTGCTTATCACTTTTAACGGCTCTATTTTCACCCACGAAACAACATTTATGACCGCTATGCGTCTGATGTTAAAAAAACTGAAAAATTCTATAATGTCGTTTATTTTCCCTTCCTACGCAGAAAGACAATCATCTGATGAAAGCGACAATTACAGACTATTACCAAATGGCTCCAACAAAGCCCAAATCTCGATAATTGACATATGGTCCATTTCCAAGAAAAGGCAAGCTGAGAAGCTGGTTCCATTGCCCATATGCCACGCAAATAGTGTGGTAGCACTGACAGGACTGCTGATCCGATCAAAGACAGAAGATCCAAAAGGCGGTATCATTGCATCCGTTGGGGATATTCTTAAGACTTTGGAGAGGTCCATCTGTGCAC tpg|BK006946.2|:214468-216301 7X167= 9S373=7X 
 tpg|BK006946.2| 567563 + tpg|BK006946.2| 566798 - INS AGTTAAGATGGAATATGTTCAGTACCTGAGAAAAGAGAAAAGGACTTTGGCAAAAAGACTTTTTGTATCTTTCAATCTTTGAAAACATATTTCCTTCACAACTGAGAAAGAGTGAATACTGAAATTGTTGTTTGTTGTTGAATAACAATACAATAACCTCTCAGTCTCAGCATCTAATCTCAACTTTACCAGCTGAAGTCCAATGTGATTGCCACCGCATTCTACTGGAGGTTCAATTGGACAAATTATGCATTCGGGAGCCTCATTCAAAAAGGAAACTGACCGATTTTCTTGGCTGCCTTCATCTTGCAAATGGGATTCTAGCAATAACCATACCGTCTCTGTCACTTTAGAATTGTTTACCAGGTGAAATAAAGGTTTATCTGCAACGATAGAAAATTTATTGTAGCGTGAAGTATCGT tpg|BK006946.2|:565940-568421 7X5=171S 10S393=7X 
 tpg|BK006946.2| 79930 + tpg|BK006946.2| 80066 - INS GGCTCGTAAAGAGTGAATTTATCGTAAATGAAGGTCTTAAAGTCACTGATGAGTTTTATTTCTTCGCTGACCGTCCATAGAAGTCTTTGCGCCAAGAAGTTACGTAAGAATGATTTCGTATATTTAACCAGAGGATCTGCACCAGGAGTCTGAAGC tpg|BK006946.2|:79604-80392 7X4=74S 74S4=7X 
 tpg|BK006946.2| 86802 + tpg|BK006946.2| 87101 - INS TAACTTTTGCTGCCATGCCACCGACGTTGAAGTTCATGAGGTGATCTGAATGGGCAATTAAGTTGTACGTCGATAGTAAATTTATGAAGCTTGTTTGGCTGGATAAAATATTGGCGAATTGTAATGTATTTTCCGGACTTTCATAATACGTGATGTTCCTATTGAAACTATCCAAAAATAAGGCAAATGTATAAAGG tpg|BK006946.2|:86394-87509 7X5=93S 93S6=7X 
 tpg|BK006946.2| 826902 + tpg|BK006946.2| 827138 - INS TTTTACTTAATCTAGGATGATGCTGTTTTTACTTCGATTTGACGTAGTAGACGTCGTGTTGGTATTTGAGATATCGGGCGTATCCACTAATAAAGGAGCCAACCCAAGTGATGCATCTACAATGTAATCATAGTCGACCCCAGAATAATTGACATTTGTCATGAAATTGTTAAAATTACCTAAATCGTTGAAATCACAGTTGTCCATTCCATGCTTTGTACTTCCAAGGATACTGCC tpg|BK006946.2|:826414-827626 16S109= 106=20S 
 tpg|BK006946.2| 114748 + tpg|BK006946.2| 115402 - INS AATGTATACTGTGTGGCCTTAGGATTTAATGCAGGTGACGGACCCATCTTTCAAACGATTTATATCAGTGGCGTCCAAATTGTTAGGTTTTGTTGGTTCAGCAGGTTTCCTGTTGTGGGTCATATGACTTTGAACCAAATGGCCGGCTGCTAGGGCAGCACATAAGGATAATTCACCTGCCAAGACGGCACAGGCAACTATTCTTG tpg|BK006946.2|:114322-115828 25S85= 97S6=7X 
 tpg|BK006946.2| 730954 + tpg|BK006946.2| 731136 - INS ATCCATCTGGCCAGAATAATGTTTTCCTATATGTACTTACCAATTATGTAGTTGAAAAATCATACACAAATAATAGCACTATAAATAACGAGCAGGATATTTATAAAAGAGTTTAACAACAGAGTTCAGGATTGAATATTCTCAGTAACTGCGTAATACATATTGTTGGGATTTACGTTTTTTGCCTTAAACCCTGTTTAATATCTGTTTAGCAAAATGAAAAGCATATGGAAACCTCTTACGC tpg|BK006946.2|:730452-731638 7X181=32S 1S1=197S 
 tpg|BK006946.2| 146648 + tpg|BK006946.2| 146672 - INS GTATAGTTCGATATGGACTTCACTACCGACAAATTGAGATCAATGGGCAGAAAATGGCAAACTTTGATCGAAGCTAATGTTACCGTTAAGACTTCCGATGATTACGTTTTGAGAATCTTTGCTATTGCCTTCACCAGAAAGCAAGCTAACCAAGTTAAGAGACACTCTTACGCTCAATCTTCCCACATCAGAGCTATCAGAAAAGTTATTTCTGAAATCTTGACCAGAGAAGTTCAAAACTCTACTTTGGCTCAATTGACCTCCAAATTGATTCCAGAAGTTATCAACAAGGAAATCGAAAATGCTACCAAGGACATCTTCCCACTACAAAAC tpg|BK006946.2|:145968-147352 7X214= 26=1X286=7X 
 tpg|BK006946.2| 54504 + tpg|BK006946.2| 54701 - INS ACTGAAATAATGATGTTGCTTCGGTTTTTTGCATGAATATAACGTGACTGTTGCGTATGCATATGTGCACGTAATTTAAAGAGAGAGTGACAGAATCTGCGCATCAGCATGGGGGCATATACAAGCATATGAGAATTTGGATAATGTATTACATCTAATTTATAAAGTTTGTAGAACAGCCTCTAATTTATTTAGTCTTTCTCCCACGCCCAATTTCGTTATTAGTTTGTCCTCCTTGCCGATTAACTCCAGCAACATTGTGGGCAACAACTCTTTGTTGTAATACCGACACCATAG tpg|BK006946.2|:53896-55309 7X204=18S 3S1=263S 
 tpg|BK006946.2| 59893 + tpg|BK006946.2| 60594 - INS ATATCCAAGGGATTTTTGAATGATTCAATTGTTTGCGAATACTCTAAAAATGTTGAACCCTGTGTTTCAGGAACACTGCCTAAAAATGATTCAAAAAAAGGAAGAAACTCGCTATCGTCTACAATGTCCTTCAATGTGATGGAGGTAAGAAATGAAGCCATTTCCTTCAATACTATTC tpg|BK006946.2|:59523-60964 10S54=32S 84S5=7X 
 tpg|BK006946.2| 866775 + tpg|BK006946.2| 867110 - INS CGAGCGTTCATAGTTCTTGCTGGTCTTTTAGTTCATTCTCTAAATGATCCAGATCTTCTTGTATGGTCCAAAGTTCGCGGTACAATGACCCTGGCATAGCCAACAGTTCAAGATGCTTACCTTCCTCTCTTACTCTTCCGTTGTCAAGGACTATGATCTTGTCTGCATCTGCAATTGTCCTCAGTCTATGTGCGATGTATACACTCGTTCTCGAACCCGAAGTAAAGTTATCTCTAATGGTT tpg|BK006946.2|:866277-867608 7X61=60S 6S1=143S 
 tpg|BK006946.2| 336120 + tpg|BK006946.2| 336343 - INS CGTATATGGACACACCCGTCATACGTAATGAGACAAAAGTGGTTGCTAACCCAACATTATCTTTGAGGTCTTCACCCGTCCAGTTACAGAGCAATGTGGATGACTCCGTGTTAAGGCAGAAACCTGATAAACCAAGGCCGATTGTTGGGGAAGAACAACTTAAACCTGATGAAGATTCGAAAAATCCTGATGAAAAAGGTCTAATGGTGCATAAAAGAAATCAATCTCTCAGCTCACCATCAGAATCAAGTTCTTCTAATCCAACGGATTTTAGCCACATCAAAAAGAGACAAAGTATGGAATCTATG tpg|BK006946.2|:335490-336973 7X245= 289=7X 
 tpg|BK006946.2| 562960 + tpg|BK006946.2| 562849 - INS GGGATTGTACACTCTAAAGGTAATACTTTAAAACTATGTCAGACGAGATTGTAACCAACAAATCTGTTACTTATGTTAACAATACTACTCCAGTCACAATTACATCATCGGAGCTGGACTTGAGATCATGTTATCAAGATGACGAAGTTGTTATAGAAGTCCATGCTGCTGCTTTGAATCCAATTGATTTTATTACTCACCAGCTTTGTAACTCCTACATATTTGGCAAGTATCCAAAGACTTATTCTAGAGATTACAGTGGTGTCATCATTAAAGCGGGAAAGGATGTCGACAATCGCTGGAAGGTTGGCGACAAAGTGAATGGTATGTACAGTCATATTTATGGTGAACGTGGTACTTTAACACAC tpg|BK006946.2|:562099-563710 15S177= 345=7X 
 tpg|BK006946.2| 693279 + tpg|BK006946.2| 693437 - INS TATCAATACAGCATTTCAGAAGCATGTCATCATTATGAATTCTTTCAGTAACTATTTTAAAAAAAAGATCAACAAAGTTCTGGTATAACTGGACGAATTCCATGTCACCGTTACACAAGACGTCGTCCAAGTTCTGGCATATACTACTAAATGCCAGTTCTATTAATTCAACAACAGATACATCATTGTTAAAATTGTTGTTGGAAAGAACTTTGTTCATAATGTACAAAAA tpg|BK006946.2|:692801-693915 7X4=112S 106S10=7X 
 tpg|BK006946.2| 150285 + tpg|BK006946.2| 150762 - INS AGATATAGAATTATTTTGAAGTTCATCAAAAGAACTTTCCTTTTTCAACGCTGGTCTTAATGGATTCTTGAATCCTGTCGATCTCGATTTTTTTTGACTGCTCTGGTCAAATGAGTTTTCAGAAATTAACTGCGGTGGTTGTATTATAC tpg|BK006946.2|:149973-151074 7X82=29S 3S1=182S 
 tpg|BK006946.2| 864439 + tpg|BK006946.2| 864605 - INS ACTGTAGTGTGTCCAATCTAATAATATGAGCCAGCGAACCTTCGAACTATGTTCTTGTAAAAACGGCTTTAGAAGATCTAGTGCATCGTCAGTGTTTCTTATTAGCGTGTAAACATCGACAGAATAATTTTCCTTTAAGTCGTTGGTCCATCCTATGGTGGCGTAATTAATCAAAGTGGTATCCAGTATTGAATTGCTT tpg|BK006946.2|:864027-865017 7X13=86S 94S6=7X 
 tpg|BK006946.2| 711269 + tpg|BK006946.2| 711626 - INS GAAATGATGAAATTCCCGCCACCACGCTTGAGAAACACGATAAAACCAATGTAACATCCGTTTTGGATGATAGATCAGAACATTTATCTAGCCACGATGTTGATAATGAGCCACACGATAATTCCATTAACATCAAAGTAAATGAAGGTGAGGAGCCCGAACATCAAGCAGTGGATATAC tpg|BK006946.2|:710895-712000 7X12=164S 90=7X 
 tpg|BK006946.2| 56439 + tpg|BK006946.2| 56539 - INS CCGAATGGGAGAATTTTGTGGGGTATTTCAATCATTGTTCCAACTTTACGTTCCTTTTTTGAATAAAGACACTTCTTATTATTAACAGGCTTTTATTTGTCAAATAAGATTCATTCAAAATTTCCATAAAGCATTACTTCTGCGATATACTACTAACGGAATTTTGGTTGCGTATTATTGTGTCTGACATTGTATGAAGG tpg|BK006946.2|:56025-56953 7X296= 100=7X 
 tpg|BK006946.2| 459705 + tpg|BK006946.2| 460157 - INS AAATTGTTTCGAAAAGACAAAAATTGTGTACTTTTGACATGATGGTCCGTGTTCTTTGATCTGCGGCAAAATGAACCTACCATGTGGCAGAATTAAATATTTGATTCAAATATAAATAAGGCGAACGACGAGAGATTAAGATATTATATACAGGTAATAC tpg|BK006946.2|:459371-460491 7X7=73S 75S5=7X 
 tpg|BK006946.2| 702546 + tpg|BK006946.2| 702826 - INS AAAACTTGTTTGTTGCCCGTTAAAACCGTTGGTGTTATGGGTGACCAAAGAACCTATGATCAAGTTATTGCTTTGAGGGCCATTGAAACTACTGATTTCATGACTGCTGACTGGTTCCCATTCGAACACAGTTTCTTGAAGAAAGTCGCCTCAAGAATTGTCAATGAAGTCGATGGGGTTGCTAGGGTCACTTACGATATAACTTCCAAACCTCCTGCAACTGTTGAATGGGAATGATTCATTTCTATTTTAACA tpg|BK006946.2|:702022-703350 13S18=1X195=15S 15S5=7X 
 tpg|BK006946.2| 176739 + tpg|BK006946.2| 176701 - INS TTGTTATTCGAAAACTAGCGACTTATTTGGATCTTTTGAGGTTAAAACATTAGAAAAATCATTTTTCTCTACACCAAGTTTCTCAAACTGGAAAAGAAAGTTGTTATTCATTTCAGATAGTGCAAAAAGATAACCGTTTTTGAAAATGTGTAATTGGTGTGAATTTTGGATTGTATCAAAG tpg|BK006946.2|:176325-177115 27S33= 91=7X 
 tpg|BK006946.2| 422342 + tpg|BK006946.2| 423004 - INS TCTATCCTCTTATGTTGGAACCGAGATATGTCTCATAATCAGACTAACTATATCTGAATTGGCTCGTTTTAATTCACGTTGTTCGTATTCACTATTCTTCATTCTAATATCATCTTTGTTTGCGATATCGCCAAACGTTTGGAAGAAGACTAGGGGCACAAGGGCGGAGTAACGT tpg|BK006946.2|:421978-423368 7X7=145S 154=7X 
 tpg|BK006946.2| 173517 + tpg|BK006946.2| 173124 - INS GAACTTTTTTAGATGAAGGAGCTATTCAAGCACCAAAGCTATCCTTCCAGGATTATTTAAGCGGTAAGGCCAAGGCTTCCCAACAGGTTCATGAAGTGCATCATAGAAAGCTTACAAGGTTTCAGGGTGAAACTTTTCTAAGAGATTGGAACTTAGTCTGTGGGCATTATAAGAGAGATGCTAAGTGTGGAGA tpg|BK006946.2|:172724-173917 7X7=16S 97=7X 
 tpg|BK006946.2| 493451 + tpg|BK006946.2| 493990 - INS CTACATGCTATATTCGTTCGTAAAACTGTTTGACATGATTTTCGAATTGGGGTTTCACTGATTCATTACCTCTTTTTAGTTCACCAAATATGAACGTGACTTGAGACGCCTCCTGCAACATGGAGCATAACTGGGTCTCTATATCATTTAATGACTTAAGACGTTCTTGTATATATGGTGGCTGCATTGTTTCGTTTTCTTGTTTCGTTTCACTCTTCGTATTGAGAACCTGCATCGTTGTTCATTTGGATTTGATAGCGTCCTTCTAATAAGCGCGCCTCTGGCTTGATGAGAAGATTTG tpg|BK006946.2|:492835-494606 7X158= 283=7X 
 tpg|BK006946.2| 19042 + tpg|BK006946.2| 19072 - INS TCAGCAAGATGCCTTGTAAGTCGTCAGATCCAACATAGTTTAATAGAGATGCAAAGGCGGCATAAACAGATGCGGTGTACATGTT tpg|BK006946.2|:18858-19256 7X12=30S 38S5=7X 
 tpg|BK006946.2| 434249 + tpg|BK006946.2| 434089 - INS GTCCATGCTGTGCCGCAGGAGAATTCGAGATGCGAATGAGCAGCAGCCATTTTGATGTTGTGAGCATCGGAACGTTTCTGCGTCCGTACACTGTCCTTTTGTTACTTAGATAATGGCTAAGGCAAGCAGTCCGGGCCACAGGAGTCAAAGGCTTTTCGCCAGCTCCTAAAC tpg|BK006946.2|:433733-434605 7X1=2I150=7S 3S1=159S 
 tpg|BK006946.2| 268712 + tpg|BK006946.2| 268106 - INS TTAGTATTAGTTCTGAAAAAAGGATTTTTAATGTGTATGCGTTCCGAACTTTAAATATAACGTCAGCGTAAAAATAATTTTTCTCCGAATGTATATCGAAATCTCAAATTGCTCTTAGAGATTTAGATTTCAACGACAGGATAAATTGGCTAGAGTTGAAAAAACTGCACAGAGTATATA tpg|BK006946.2|:267732-269086 7X5=247S 158=7X 
 tpg|BK006946.2| 717843 + tpg|BK006946.2| 717836 - INS AATAAAACAAAAAAGAAGAAAAAGCTATGCATATTCCTATCACAGTTAACGCTTGCTTCCGTTCTTTTTTCTATATCATCGTTTCCATCATGTTTTTCTTTAAATTGAATACTTTCCTATGCTCTTAATGAGTTGCGATTGTGCATATACTGTATTTCAAAATCCTTTGTAT tpg|BK006946.2|:717478-718201 7X45=41S 6S1=169S 
 tpg|BK006946.2| 370110 + tpg|BK006946.2| 369670 - INS GCGTATAGCTCTTACAATTTTCATAACTCTCTTGGCTTCGTTTTTGGATGGAACAAATCTTCTTTTTGGCTCCGGAACAGCAGTTAATGGCATCACTTCTTCGTGTCTCGTGAACCAATCGATTAACGGTTCGTATGGATTTATGCTATCATCAGTTTGTTCGTTCCTTTGGATTTTGGAAATAAGTTCTAATTCCTCTTTGGTTAAGTTCAAACTTGAACCGGAATTCTTGTCCAGTAAACCAGTCCAGCCTTCAGGTAGCTCGATAGAATCCAACAGTTGATCTAAAGC tpg|BK006946.2|:369074-370706 7X6=150S 146=7X 
 tpg|BK006946.2| 503094 + tpg|BK006946.2| 503011 - INS GTGATTCTCTTATTATGAGGACTATATTGCATGAGAACTGGATGCGATGCAAGTACTTCTGGTACAAACATGTAAATACTAGTGATTATATTACAGTAATTTTGTCAAAACACAGTGGCACAAAGTCATTTGATAATGTGATAGGATAACGAAACATATAAAGCGGAAGGACAAAAAAAAAGTAGTGATATTATGTAGAAATACCGATTCCATTATGAGGACTCTTATATCTTCGAGAGGAACTTCTATTATATTCTGTATACACAACATTATAGCCTTTGATCAACAATGGAGTTCACAATTATCAAAATATTCGCACAATATTCACGTAGAATAGTGGATGACAGAGTATATAAACAAAGAAAGAAGCACTCAGGATTTTCTATAAATAGTGAAGTTTTCTATGGACGCCAAAAAATCTTAAGGGTATCTTGAGTG tpg|BK006946.2|:502121-503984 7X3=174S 7S61=1X356=7X 
 tpg|BK006946.2| 707657 + tpg|BK006946.2| 707695 - INS ATTCCAGTGAAGGACAGAATTATTCAGAGGGAGTAGAAATGGAATTAGAAGACGACATTGATGTGGAAAGCGATGCTGAAAAAGATGAAAGTCAGGGTGCAGAAGGAACAGAACATTCGGTAGATTTTTCAAAATACATGCAGCCTAGAACAGATAATACTAAGATCCCCGTTATCGAAAAATATGAATCTGATGAGCACAAAGTCCATCAAAGATATTCAGAAGACGGTGCATTTGATTTCGGTTCAGTAAATATTTCAG tpg|BK006946.2|:707121-708231 7X130= 196S4=7X 
 tpg|BK006946.2| 467409 + tpg|BK006946.2| 467549 - INS AAAATGGGAAGATTTTCCAAGACAATTTGCAAAATGTCGTCGATGCAAAAGAACGAAATATTGCTCACGAAAGTGTCAATTAAAAGCATGGGGATATCATAGGTATTGGTGTCACGAAGTTGGATCAAGTCATATGAGATCCACGAATACTACCACAGGTGTCAATACCCCAAATGAGCCTAGTTCTTTAAATGCCACCGCTACTACAGCAGCTGATGTTTCGAATTCTACCAGTAGGTTCACTCCTAATATATCCACCAGCGTAC tpg|BK006946.2|:466863-468095 7X236=1X6=6S 9S1=258S 
 tpg|BK006946.2| 33547 + tpg|BK006946.2| 34176 - INS TAAAGAGAGGATGCCG tpg|BK006946.2|:33501-34222 7X6=2S 8=7X 
 tpg|BK006946.2| 486715 + tpg|BK006946.2| 486816 - INS GTCTAGACGAGTTCATAAATTTTGACCCAGAAGTTGAAAGACAACAGACTGAATTACGTCATAAGCGTACAGGCGGTAAGCACTGAATTTCAAAAACATTTATTTCAAAAGCATTTTCAGTAAAAAATGCAGACTTTATTATTATTTAATCGTGCTTCTTATATATGACATTCTACCAAATCG tpg|BK006946.2|:486335-487196 7X5=86S 89S3=7X 
 tpg|BK006946.2| 749591 + tpg|BK006946.2| 749866 - INS ATGCGCCAAAATAGTTTCTACCCTGTTTCTTGGACCTTGAATGGTGATTAGGGATTATTTTTCCGTAAACGTCGCCTTTTAAATTCGTTATATCCCAATTCAAGCCGGCAATTTTCAGATCAGGATATCCCGTAGGTAATCCAATGTCTTTCATCTTCATACACCATGGTGGTAGTT tpg|BK006946.2|:749223-750234 7X93=39S 1S1=35S 
 tpg|BK006946.2| 321233 + tpg|BK006946.2| 321374 - INS GAGTATATATATACAACTATCAGAAGA tpg|BK006946.2|:321165-321442 7X3=10S 14=7X 
 tpg|BK006946.2| 846043 + tpg|BK006946.2| 846250 - INS TTCATCAATGCAGCATGCCACTCACGGAAGTCTTGGAAAGCAAGGCATACTGGCATAAAAATTGTGCAGCAAATAGGTATACTTTTGGGAATAGGTGTCTTGAATCATCTTACTGGGCTGATGAGTTGTATCAAAGAC tpg|BK006946.2|:845753-846540 7X25=44S 2S1=165S 
 tpg|BK006946.2| 780952 + tpg|BK006946.2| 780740 - INS GCAATGCAATGACCATCAGTCTATGCTAATATTTGAAAAGTCCTTCGAATTGATTGGTGTTGACAAAATACCTAGAAATGCACAAATGAAACGAACCGTCTATGCTAATATCATTATCTCTCTGGATTTTTTCCAAGATTACTTTTAAATTCTCGAAATTGTTAGTAGAGACGTACGCTTGAACCACTGACATATATAGCTCTTTTCGTGTTGAAATATTATTATTAAGTCTGGTAATAAATTTATCAACTCTTTCCATCAATATTGAGTCATCAATGCTTTTTGTTCTGTCTCCTTTGATGCAATACAGAGA tpg|BK006946.2|:780100-781592 7X7=10S 7S287=7X 
 tpg|BK006946.2| 216220 + tpg|BK006946.2| 216404 - INS GCCCAAGCGATAACATCACAGTTATACGTTCAAGATGTCACGCATGCCATCTAGTTTCGATGTTACGGAGAGGGATTTGGATGATATGACCTTTGGCGAAAGGATTATATACCATTGTAAGAAACAGCCATTGGTACCCATTGGGTGCTTGCTGACTACAGGAG tpg|BK006946.2|:215878-216746 7X63= 82=7X 
 tpg|BK006946.2| 895049 + tpg|BK006946.2| 895593 - INS GGAATAGAGGTGTCTCTCGTGGTTAAGGGAACATATACTGATTGTGTATAACCCTCTTTTAAAGGCCCCTTCATAAACAAGTCTGTGAACGATGACGCTATACGAGTATAGTAGCCATACTGCGAGTCCAATCCGGTGAAATCACCGTAAGCTTCCTGAGGAGATACAATTTTCCTCGTTATTGTGTCGATGGTGACCCTTGCGTTTATCGGCACCAGCTGACTTTGTAGAGCCAGTGCTTTGCTTTTCCCTATATTAATATATTTGGTTTGCTTGAATAC tpg|BK006946.2|:894473-896169 7X231=23S 4S1=176S 
 tpg|BK006946.2| 121389 + tpg|BK006946.2| 121320 - INS CCAATAATTTCATCCTCATCTGGGGTCAAGTCGTAGTCTTCACTGTCATAGATGTCAGCGTCTTCATCTTCGTCTTCACCTTCGACTCCCATTGGAGTATCAAATGGATGCTTAACATAGTTACCGCTCAAGGAGATAGCGTAAGAACCAGTGACAATGAATTGGACTTCTTCTTCTGGAGTAATG tpg|BK006946.2|:120934-121775 7X4=89S 89S4=7X 
 tpg|BK006946.2| 477770 + tpg|BK006946.2| 478428 - INS CCTCTTTCTTGATGCCGAGCACTTCAACCAATTTTGTGCTATCAAATTTCTTGTGCGTGTAAGGACTTATTTTGTTTTTCAATGAGTCAGGAAGCTCTGGGATTTCAAATTCCCTGGAATCATTGATCATCAGTTGGTGAATCCATTCCAGTAGCACCTGTTGTTGCCTGTAGACAAAAACCGTGGGTATTCTAAGAGGATCCTTTTTGTTTTCCTCTTGGTCTTTATTTAAAGAGGGAAGTGGGAGAGTGGTGTCTGTTGTTACTTCGCCTATGGGTTGATAGTAGTTGCCTAACGGAATCTCTGGTAGCTCATCTGTAT tpg|BK006946.2|:477114-479084 7X18= 161=7X 
 tpg|BK006946.2| 648840 + tpg|BK006946.2| 648898 - INS ACTCTATGATTTCAGAACTAGAAAGGCTTATTGAAGAAATAAAAACTGCAAACAAAAATGGTACGTTATTCGAATATTCTAATTCTAAAAATAATCCTTTGGGAGCCGGCTGGTCAGGATTTAAAAAGGTTTTTAAATAGTTAAACTGTGTATATCAGCTACTGCTCCCCTTGAATGATAC tpg|BK006946.2|:648464-649274 14S127=24S 19S4=7X 
 tpg|BK006946.2| 311402 + tpg|BK006946.2| 311876 - INS GTCGTATCACTTATGCTAGTTCTTCTCAAAAATATAAGTTCCTCTTGCAAGAATATGAAGGTAATTTCACTTTATCGCGCAAGTGCATATTTCTGAGTTTACTATGTGCTTCGTCTGAAACCTCTCATTATCTACTTAATATCGGCTATTCATCTCACGTATTCACGTAATATTTGATTTTTGTACTACTATTTCTCTCTGTCATACGTGCATGATACATTTCCTTGTTCAAATTAAAAGAGTCACCGTCAGC tpg|BK006946.2|:310882-312396 7X21= 238=7X 
 tpg|BK006946.2| 404442 + tpg|BK006946.2| 404665 - INS GTATATTCTAAAGGGTTTGAAAAGACAATATTTACGAGATATTAGTAACATCAGTAAAGATGCTTGTGAGTACAAGTTACGGAAGGCGGAGCTAATGAATAATGAGTCAATCTTAAAAAACATTCCACAGGGTACAAATCAAGAGAATACAATAT tpg|BK006946.2|:404118-404989 17S12=55S 73S5=7X 
 tpg|BK006946.2| 177501 + tpg|BK006946.2| 177572 - INS TTACCAGAATCGGAAGTTAGCGCTAGAAAAGTGGGCCAGTTGGAAGCTTTTGCCCTTGACCCTGAATGCGGCAGATCCAGCGACTTCATCGAGGTTATCGTCGCAAACAGGTTTTGAAACTTGGCAATAAGCTTTAGTTCCCCATCTGCAGTATCATAAAGTTCTAAATGCGTCTCAGTAGCTA tpg|BK006946.2|:177119-177954 7X116=22S 1S1=213S 
 tpg|BK006946.2| 691492 + tpg|BK006946.2| 691515 - INS AGATTTCACTGATTGAGAACCCCGAAAAGAGCCATCTCTTTTCATATTATTTGGAATATTCTTTTCATTCATAGTTTTTTTCAAATCGCTAACTTTTGGTGCGGTGGCTCTCATTGTTTTCCATGATCTTGCGTCCTCAGCAACAAACCTATAGATA tpg|BK006946.2|:691164-691843 7X4=74S 75S4=7X 
 tpg|BK006946.2| 784746 + tpg|BK006946.2| 784697 - INS CAAACTTTTTTGTGAATATAAGAGCGGTCACACTGGTGTTCCTGTTATATTCCCAGTCTGCAGTTTGAATAAAGTTCTTATTCAAATAAAAAGAAGCCTTTTCTCTTATTTCAGAATCATCGTCCCATAAGAAGTTGTACAGTTGTAATAGTATTCTGGAGTTCTTACAACTTTCTGGATAAGCAGTTAAACAT tpg|BK006946.2|:784295-785148 7X91=54S 2S1=251S 
 tpg|BK006946.2| 807069 + tpg|BK006946.2| 807142 - INS GTTCTATTGAAAAAATATTGCGACTGCCTGCCTGAATTCAGCTTGAATGACCCAAATCTTAGTGCTTTGCATTCTAATCCCAGTTCAAGGAAAGTTTTTTGATATTCCTCTAAACTTGTAGTAGATGCAGACATTATTGGATTATGTTTTATTATTCTTGATGGCTCTAGGTCTCGACTATTTTGCGTGACACTTCCTTAGTTCTTAATCTATATAAAAGAGCCTGTGA tpg|BK006946.2|:806597-807614 12S13=1X181=14S 11S4=7X 
 tpg|BK006946.2| 735193 + tpg|BK006946.2| 735326 - INS ACATACAAACCATCCACTTTTGAAGTGGATCTGGACCGGAGAGATACGACGGGCGATTTTTCTGAAAATATTAGAACAGTTTTTTACAGTTACAAAACATTCTTCAACTACATGAACTCAAATGGTACATCAGACGCAATGAGCGAGTCTTCAGAGG tpg|BK006946.2|:734865-735654 7X6=3S 79=7X 
 tpg|BK006946.2| 748381 + tpg|BK006946.2| 748723 - INS TGCATACCCTGGCCCTAATCGCTAAATCTTGAATCTCTGGTAATTTTGGAGGCCATTTTGTTGCCTTGACGATATCACCAGCCTTTGTTGGGTCATAGCTATCTTCTCCTTCGTCTTCTTCTTCATCTTCCTTTTCATTTAAATTTTCGTACACATTTACATCTATTTTCTCTCGCTTTTCCCTTTTAACTTGTTCTAGCTTCTCTAACTTTTCCATATCAGCTTTACTGATTTCTTGCAATATAGGTTGCTTT tpg|BK006946.2|:747859-749245 10S211=16S 19S5=7X 
 tpg|BK006946.2| 108053 + tpg|BK006946.2| 108211 - INS AACAAGATTGTCATCAAGAACATTGTATTGCGGTGCTAGAATTCTTGGCGATACACCAGTCTGGCCCGTATCTCTGTTGTTTGCTCATGCCTTACAATCTAGGGCTATTTACAATATCAACCACAGGAAATCTGTAAACAGTGTATAGACT tpg|BK006946.2|:107737-108527 7X132= 6S1=7X 
 tpg|BK006946.2| 556985 + tpg|BK006946.2| 556467 - INS GAATACAATACTAAACATGCAAAAGAAATAATGAAGATAAAAACAATCGACACACTTATAGTTCTAGCCCCAACAGCACAAAAGCGGAAAAAATCAAAATCAAGAACAGGCCAATGAGCGTTGTCTTATATAACACAACCTCTTTTATATATACACCCAAGAAGGAGAATGAAAATAGAAACACCACACGCTTCGAGACAACGGAAAGAAAGCATAAGGAGTGGCCCATGTGTGCCAAAACTCTTCTCATTGCCGAGCCATGTATTACCATCCCGATGGTGATGGTTGTGAATGCAAATACCGCTGAGGCCAGAGTAATGCCATAGCGAGGACCAGGGCATCTCGAGCATCGTGGAG tpg|BK006946.2|:555739-557713 7X5=159S 179=7X 
 tpg|BK006946.2| 729127 + tpg|BK006946.2| 728881 - INS ACTCTGCCATGCCGATTCTGATCTTTTTCAACTGAGCCCTATTTTGTTCAATTCTGGAATCAGAGAGATGACCAACGTAGATGACACCACGCAAGCCAACATCAGGAATTTCAACAATAACAGAATCTTTGGTTTTTTCGATAACATGGACAGTAATGATTGTTC tpg|BK006946.2|:728537-729471 7X3=149S 11=1X143=7X 
 tpg|BK006946.2| 421425 + tpg|BK006946.2| 421645 - INS GTTCATTGATTCAGGATAAATATATAAAGAAAAAGCCACTATCCCCAGAAATTTTGCTGTTGATGAAGGCTACGATGCTGTGAATTCAGATTATAGGAGAAATTCACCTCGAGGACTTGAAATCCACATTAAGGAATCGATATTTTT tpg|BK006946.2|:421117-421953 7X6=67S 67S7=7X 
 tpg|BK006946.2| 313406 + tpg|BK006946.2| 313434 - INS TTCTATTTCAGAACCTGTTACAGACAGACGGCGTGCTGGAACGCGTTAAGTCAAGCGGTGAACATGTGTAATGGGATGAGTCTATATTTAAACAAATTTCCTGAGATCCATTCCACTTATGATGAATCAAAAGCATGGCATTGTTTCTGGTGTTGTTTTATAATGGATAAGTTGATAAGTTTTCAAATTGGTCGATTCTACCAACTATCATTACCCGCGAGCGAGATG tpg|BK006946.2|:312936-313904 7X180=19S 2S1=246S 
 tpg|BK006946.2| 706604 + tpg|BK006946.2| 706920 - INS AGGGATACCCTGTT tpg|BK006946.2|:706562-706962 7X3=4S 1S6=7X 
 tpg|BK006946.2| 501405 + tpg|BK006946.2| 500814 - INS GTCTTAGCTTCAATTTTAGAATATTTTCGTTTGCTTCCGGGGTGACCGCACTTTGTTCTTCCAGCTCAGGTTCAATTACTTTTGCTTTTATTTTGGAACCGTTCGGTGTGGATATTATTTCACTATCTTTGAGGTACAATTTCATCTTTTCGTCCAATTC tpg|BK006946.2|:500480-501739 23S18=1X211= 80=7X 
 tpg|BK006946.2| 223896 + tpg|BK006946.2| 223730 - INS TCACACCATAGTATACTAAGGACCTTTTCCAGTTAGGATAGCAAAGGTGTCAGAATTACCATAGCCCAGGCATCAACCAGTTTCCGCGCAAGAATTCTCCTCCTCCCGGAACAAGAGGCCTGCGGAGACGAGTTCTTTGCCTCTGAAAGGCGAATCTCTGGAAGGA tpg|BK006946.2|:223384-224242 9S164= 146=7X 
 tpg|BK006946.2| 737751 + tpg|BK006946.2| 738329 - INS CCCCCATTGTACTACCGTT tpg|BK006946.2|:737699-738381 7X6=3S 7S3=7X 
 tpg|BK006946.2| 586439 + tpg|BK006946.2| 586505 - INS GTATAAAGAGGCACCGTCTTTGTAGCTGGCCAGATAGCTTGCTTACCTATTTTCTTGCTAGTTTAAATTCGACCGGAATAGAAATTTGGTTACAAGAACGCTATTGCGCACCAGATGCAAATTTTTTTTTTATTTTATATAGTGTCACTGGCACCCCTCCATTACATTGTCTAATTTAAAATAACTAAACTGATATAC tpg|BK006946.2|:586029-586915 14S14=1X105=21S 46S4=7X 
 tpg|BK006946.2| 481014 + tpg|BK006946.2| 481336 - INS TGCAACCGATAAACCATTATAAATCTTCGCGGTTATCTGGCATTGTTATTAACCAAAAAAATGCCGGCCTATTACAAGCTACTGTTCAATAAATATTGTTGTAATGAAGACGGTCCAACTGTACAAATACAGCAAACTGTCATATATAAGGAGTCTTATGTGACAGCACTTGCGTTA tpg|BK006946.2|:480646-481704 7X5=83S 84S5=7X 
 tpg|BK006946.2| 253383 + tpg|BK006946.2| 253607 - INS ACCATGAAGAGTAGGAGGGTGGCAACTGATGGATGCGTAAGGTCTTAAGAGATACATTTGCTTAATAGTCTTCCGTTTACCGATTAAGCACAGTACCTTTACGTTATATATAGGATTGGTGTTTAGCTTTTTTTCCTGAGCCCCTGGTTGACTTG tpg|BK006946.2|:253059-253931 186S36= 78=7X 
 tpg|BK006946.2| 544500 + tpg|BK006946.2| 545239 - INS TGTTTATATTATAACGATGGTATAATGCCTACTGTGGGTTTTCAAATACATAGTCTGATGATAAAAGATGTGACAATATCTCTATGGGACATTGGGGGGCAACGCACATTAAGGCCATTTTGGGATAACTATTTTGATAAGACACAAGCGATGATATGGTGTATAGA tpg|BK006946.2|:544152-545587 15S35= 147=7X 
 tpg|BK006946.2| 815549 + tpg|BK006946.2| 815981 - INS AAACTACTGAACAACCGTTACCTGTGTGCGATATTGAATCCTCAGATAATGCGTGCTTTGAGTGTTGTTTTAGGGTACTGACCTGTTTTTTAAAAATGTTGGATAAGTTGTGAACACTAACTTTCAAGTTGCAAATGCTTTCGATATCGTTAAACAGCTGTGAAG tpg|BK006946.2|:815205-816325 14S5=1X69= 83=7X 
 tpg|BK006946.2| 908173 + tpg|BK006946.2| 908347 - INS AGAAGGAGTCTAGCGTAGTGAGTTCAGAAGCTCCATCGTCAACATCTAGCTCAGTGAGTTCAGAAGCTCCATCGTCAACAACATCTAGCTCAGTGAGTTCAGAAGCTCCATCGTCAACGTCTAGCTCAGTAAGTTCAGAAGCTCCATCGGCAACGTCTAGCGTAATTAGTTCAGAAGCTTCATGGGCAACGTCTAGCTCAGTGAGCTCGGAAGCTCCATTGGCAACGTCTAGCGTAGTGAGTTCAGAAGCTCCATCGTCAACATCTAGCTCAGTGAGTTCCGAAATTTCGTCAACAACATCTAGCTCAGTAAGTTCAGAAGCTCCATTGGCAACGTCTAGCGTAGTGAGTTCAGAAGCTCCATCGTCAACATCTAGCTCAGTGAGTTCCGAAATTTCGTCAACAACATCTAGCTCAGTAAGTTCGGAAGCTCCATTGGCAACGTCTAGCGTAGTGAGTTCAGAAGCTCCATCGTCAACATCTAGCTCAGTGAGTTCAGAAGCTCCATCGTCAACAACATCTAGCTC tpg|BK006946.2|:907107-909413 7X4=295S 91=36D288=3I13=7X 
 tpg|BK006946.2| 73169 + tpg|BK006946.2| 72992 - INS ACCAAGTTCCACAC tpg|BK006946.2|:72950-73211 7X4=3S 3S4=7X 
 tpg|BK006946.2| 194416 + tpg|BK006946.2| 194420 - INS CAATTGGTGACGGTTATGGTTGGTCTCAAGTAAATGACAACGGGTTTGGACTGGCATACATGTTGAATAACGAGTGGCTGCATATCAATATTGTCAAC tpg|BK006946.2|:194206-194630 14S35=31S 20S5=7X 
 tpg|BK006946.2| 12942 + tpg|BK006946.2| 13474 - INS CGATATTTAGCAAGCATTTCTAGTTCTTTATGTGGTGAATAAGTAATGTGTGTGGGAACTATGGCTACTGGATGACTATATTCGGCATTAGTATTTAATAAGGGTACGACTCTGAAGTATCAGAGTTGCATCATTTCAGACACACTGGAGGGATCCTGTTATATATTTTGAAATAAATAATGTACAATTTGACGGGTGTACAC tpg|BK006946.2|:12522-13894 7X54=1X8=38S 1S1=213S 
 tpg|BK006946.2| 557261 + tpg|BK006946.2| 557137 - INS AGCATAACGTAATGAAAAGGCTAAATATTATAATGACTTGCACTTCGTATCAAGATATGCGAGAGATCATCATAAACGAAATAATATCCACAGTTTGGGTTTCATATTCTTATATATATATACGTGCGTATATGCATATATGTATGTTTACTATACATCAACATCAGCATCAAAATTAACATTAATTAGCTTCTTGCATGTGCTCTTTAGCTT tpg|BK006946.2|:556697-557701 7X106= 107=7X 
 tpg|BK006946.2| 327264 + tpg|BK006946.2| 327879 - INS AAACTGCAGTAACTTCAAGGATCGTTATAACCCTCAGCTTAGCGAATTGTACGCGCAACCAAAAAATAACAAAGATTTATCTGGAGCACAGTTGAAGAGAAAAGAAAAGATTGAGCTATTCCAGCGCAATAAAGAAATTAGCACAAAACTGCACTGCTTGGAGTTGGAATTAAAAAACAACGACGAGGACCACGACCATGATGAATTACTAAGAGAACTATATTTGATGAGGTTACATCACTTTAGTCTTGATACGATTAACAACAT tpg|BK006946.2|:326716-328427 7X7=13S 251=7X 
 tpg|BK006946.2| 768953 + tpg|BK006946.2| 769025 - INS CAATACTGTTCTTAGACAATTATCCAACCATCGCCATTAAATGATAAAAAAATAAATTGACTGCTTAATTTTGCTGATACAATGCACTATATTATCGGCTGATGTAATGGTATTGTTATTCAACCTCCTCTCGGCATTGCAACATACTAATAGCCACCCTAGGGTGTCATTAGCATGCCTATAC tpg|BK006946.2|:768571-769407 7X5=87S 87S5=7X 
 tpg|BK006946.2| 898399 + tpg|BK006946.2| 897935 - INS ATTTCATAATTCATTTTTTTGTTCAATAACAAGAACCAAACATAAAAAAAAATACTTTAAGAATAAACAAGACTGATGAAGCATAGATCATATTATTAGAGCGCGTAAGGTATGTAGAGCACAGATTGGTCCTTCGAGTGTGATTATATAATTTTATATACGCTCCTTAATTTAAAAGCGGCTTAGATAGATTTTTTATACTTTGCTGTTGGAAAATTCCTGCTGAAGCAAAAGAATTTGCAATTCGTTCTTAGCCTTTAACC tpg|BK006946.2|:897395-898939 13S125= 132=7X 
 tpg|BK006946.2| 805033 + tpg|BK006946.2| 805299 - INS TTAGAGCATCTTCCGTC tpg|BK006946.2|:804985-805347 7X1= 13S3=7X 
 tpg|BK006946.2| 440224 + tpg|BK006946.2| 440050 - INS TGTAAAAGGCAGTTATTCGGCCCAAGGATCAGTTGAAAAC tpg|BK006946.2|:439956-440318 7X10=10S 13S7=7X 
 tpg|BK006946.2| 774965 + tpg|BK006946.2| 775249 - INS GGTGTGGCTCGGTGTGCAATCGGGTGTAGAAA tpg|BK006946.2|:774887-775327 7X6=10S 1S15=7X 
 tpg|BK006947.3| 732329 + tpg|BK006947.3| 732364 - INS CCGTGTGGTCTTACTATAACCCACTTCATCAATCATGTGCGTAGCAGAGTCAATGCCAACAAATGCCCAGATCGGATTGACCAAACCGACAACAAACGCCATTCCAGACGAATTCCAGCCTGTTTGATTATCAAAGCTCCCAAATATATTAGAAGCTTTGGGCCATGGGTCTACGGTGTTGTCAGATCTTGAAACAATACAAATAATGAAAGTCATGGCGAAAGACAATAGAGACGTATAGAGCCCAAACTGAGAGATATAGGGCAACGGAGTTGAATAAATGTTGAAA tpg|BK006947.3|:731737-732956 30S292= 271=7X 
 tpg|BK006947.3| 662966 + tpg|BK006947.3| 662763 - INS TTATAGCTGCCGTGGGCAGCACATTAGGTCCCAATTCAACATATATAATATAATGCATGTCGACACCGCTAGGCTGCATCCTTTGGCTGGTCTAGACAAGGGTGTGGAGTATTTAGATCTGGAAGAAGAACAACTATCCTCGTTAGAAGGCTCACAGGGTCTGATCCCTTCCCGTGGGTGGACCGATGACCTATGTTACGGTACCGGTGCCGTCTACCTGCTGGGACTTGGTATCGGAGGGTTTTCTGGTATGATGCAGGGTCTGCAGAATATTCCGCCCAATAGTCCCGGAAAATTGCAATTGAACAC tpg|BK006947.3|:662131-663598 7X502= 23S258=7X 
 tpg|BK006936.2| 255162 + tpg|BK006936.2| 254787 - INS CCAACAAATACTACCTTTTATCTTGCTCTTCCTGCTCTCAGGTATTAATGCCGAATTGTTTCATCTTGTCTGTGTAGAAGACCACACACGAAAATCCTGTGATTTTACATTTTACTTATCGTTAATCGAATGTATATCTATTTAATCTGCTTTTCTTGTCTAATAAATATATATGTAAAGTACGCTTTTTGTTGAAATTTTTTAAACCTTTGTTTATTTTTTTTTCTTCATTCCGTAACTCTTCTACCTTCTTTATTTACTTTCTAAAATCCAAATACAAAACATAAAAATAAATAAACACAGAGTAAATTCCCAAATTATTCCATCATTAAAAGATACGAGGCGCGTGTAAGTTACAGGCAAGCGATCCGTCAGGTGGCACTTTTCGGGGAAATGTGCGCGGAACCCCTATTTGTTTATTTTTCTAAATACATTCAAATATGTATCCGCTCATGAGACAATAACCCTGATAAATGCTTCAATAATATTGAAAAAGGAAGAGTATGAGTATTCAACATTTCCGTGTCGCCCTTATTCCCTTTTTTGCGGCATTTTGCCTTCCTGTTTTTGCTCACCCAGAAACGCTGGTGAAAGTAAAAGATGCTGAAGATCAGTTGGGTGCACGAGTGGGTTACATCGAACTGGATCTCAACAGCGGTAAGATCCTTGAGAGTTTTCGCCCCGAAGAACGTTTTCCAATGATGAGCACTTTTAAAGTTCTGCTATGTGGCGCGGTATTATCCCGTATTGACGCCGGGCAAGAGCAACTCGGTCGCCGCATACACTATTCTCAGAATGACTTGGTTGAGTACTCACCAGTCACAGAAAAGCATCTTACGGATGGCATGACAGTAAGAGAATTATGCAGTGCTGCCATAACCATGAGTGATAACAC tpg|BK006936.2|:252983-256966 7X22=1X18=1X64=1X13=1X213=1X24=1X10=77S 554S13=459S 
 tpg|BK006947.3| 743992 + tpg|BK006947.3| 744656 - INS AACTGGGTATATGTTACATTGATTTATGCTTCAAGGCTTCGGATGCTCCAATCATAAAAGCTTGTCCCAGCAATGAAACAAACAATGCAAAGATGGACAGAAAAACTTGACCGCTGTACAGCGAATCTTTTTTCTTTACCTCAACGGTCTCACTTCCAGTTGTATCTGACTCTTCTAATCCGCCATCTTTGGCTCTGCCGCAGGAGCACCCGACGTTTATTAACTTTGGAGCGAAATAGCTTCCAGTCACACCAAGTATAGATGCGACCATAAACGCTATGCCTTGAAACTTGGTGTCCCAGTTAACGTGGAGCGTCAGGAATAGTGGCATAAAATAAACTACTTCGCTCATAATAAATGACGATAGGAACATGCTCCATAGTAAAATCAAGCAGGAGA tpg|BK006947.3|:743180-745468 7X337= 4S383=7X 
 tpg|BK006947.3| 177080 + tpg|BK006947.3| 177634 - INS GTCTGAAATTCGTTTCAATCATGAACTCTGAAGATGGTATTCAAACTGTTGATGAATTAAGGGACCAACAAAGGAAGATGAATGATTCTTTACGTGAACTGAGGAAAACCATTTCAGATTTGCAAATGGAAAAAGATGAAAAGGTGAGAGAAAATTCAAGAATGATTAACTTGATTAAAGAAAAGGAATTAACAGTTTCTGAAATTGAATCATCTTTAACACAGAAACAAAATATTGATGATTCTATAAGGTCAAAAAGGGAAAACATCAACGATATCGATTCTAGAGTAAAGGAGTTAGAAGCACGTATTATTTCATTAAAAAACAAAAAGGATGAAGCGCAAAGTGTTCTAGACAAAGTAAAAAATGAACGTGATATTCAAGTA tpg|BK006947.3|:176294-178420 7X333= 4S358=7X 
 tpg|BK006947.3| 548270 + tpg|BK006947.3| 548790 - INS GAGCACTTGGATGACAGAACATGCAGTGAAAGCAGTAGTAGAAACGAAAGCCCCGTAAGAACCATCACAAAGGATAATTCTGTAGGCAAGATTTTAAATAGTACTTGAGTGATCATTATTTTCTTTTTGATGTTCCCCCTACGTATGTATACACCCATATATTATATAGATACCCGCCGCATACCAACATAAAAAAGGTAACAAATATTTGAGATATAGAGCATCGCTACATTATGGGCAAGATGCGTCTTTGTGAGACGATTTTAAACAGAAGTTGTTCATCTCTCAGTGATCAATACCTATCAACATGTCAAATTCATCAGTGGAAAAATTTAAAATTTCGAATACCTGATC tpg|BK006947.3|:547548-549512 7X2=2X326=12S 4S1=233S 
 tpg|BK006947.3| 264512 + tpg|BK006947.3| 264809 - INS GTCCCATGCTTCTAACACAACCCATGTCTTCAATTAACATTTTCCTTAACCACTGCGTCTCTTGGCGCTGTAATTCCAATTCTCTTTCTAATTGCACAATTCTTTGGCCTTTTTCAGAAATGATTGCGTCATAAGCTTCTTTCAATGGGCGTATCACGGCTTCTGTATCTATAGGTCCCATGCTGTTTGAAGGATTTAAATCAACTTTCATTTGGGTGTTATTCGCGTTTAAATTAGTGTCCGGACCATCATTTATTAACGCACCCTCTGCTGCAGTTGTCATCGGCCTCTGCCTCTTACTCGTATTTGTCAGTTGCAAAAGTTCTTCCACCGCTTCGTCATCCAGCGTATTAACATCTAACGATCCCAGTGACCTTCGTTTCCACGAATGGGATCCATTATTGGACATTGTATTATAGCCCATGGTATTACTGGAAGCATTGGGGTTCAGATCTGCATGACTCAAACCAAATTCAAATCCTCCTGAGCCAGGACTGGTTGGCTGTGTATAATAT tpg|BK006947.3|:263468-265853 7X447= 499=7X 
 tpg|BK006947.3| 351962 + tpg|BK006947.3| 351455 - INS CCGCATACACATACTAAGCATAGGTACACATACACCCCTCTTTACATATTCTCAATACCTGACTGACATAGTATGCGCTACATAGTTTTGTCCTATTTTTTTTACACCGCGATTTGAAGTCTAAAGCCAGAGAATGAGGAAAAACGAAACAAACTGAGATCATTTGTATAAGGGGAGTCACTGTACAGCTGCCAATACCAATTTTCCTTCTGCCAAATCAAAAAAGTATCCGCATACACATACACCCCTCCCTCTACAATCTTAATTATTTACTGATTCCTTTCGTATTTGTCCAGTATGAGCAATACTAAGCATACCACTTCTCATCACATGGAACTCAAAAGGATCATTATCCTTACACTTTTATTCATACTCATAATGTTGATATTTCGAAACTCAGTGTCCTTCAAAATGACATTTCAAGAACTACTGCCACGATTTTACAAAAAGAATTCAAACTCAGTTAGTAATAATAACAGGCCCTCATCTATTTTCTCGGAAAACTTGGTGGATTTTGATGATGTTAACATGGTCGATAAGACCAGACTGTTTATTTTTTTATTTTTCAGTTTCATCATTACTATAC tpg|BK006947.3|:350269-353148 7X5=181S 11S548=7X 
 tpg|BK006947.3| 486572 + tpg|BK006947.3| 487341 - INS GGAAGTTTTCTAACGTACGACGGCGATGGTGATGATTTTGCATGTTGCAAATGGGGTTCAAGATGTACTCTTGATGTGCTAGCGAGCTTGTGGTGGAGTTCGACGCCGACCTAGACGTTGGTATGACGTTATCTAGCGGAGAGGAAACATTATTGGAGTTCTTCCTCAACGATGGAGTTCTAACCTCGCTACCAGAGATAGGTATC tpg|BK006947.3|:486146-487767 7X1=2I16=84S 3S1=196S 
 tpg|BK006947.3| 731306 + tpg|BK006947.3| 731589 - INS AGAAGAACAACTAAGGACTGTTTTTCTTTCAACAGCATCTTAGATGCATGTAGGGAAAACAACGATGCTGATAATGCAGAAAACTACTGCATACACTACTGAGGTGTAATTCATGTTTCCTGCAGTAACCGGTAGTGTATATGGGAAAGATAAAAATACCAGGCAGAACAAGGTCCATAGAATACATATAATATGAGGAATCATAGACATACGACGACGGTTAGGCCTGCTGACACAATTTACGTCACTCTCGATTCTATGAATGAATTTTTCCTTTTTAATAACGAACAGGAATATAAAAGAAGGAACTGCGTACGACATTAGTAACAGGGTGATGCATGCAGTGATAATTGCGTTGAAAGCGGTACTAGATCCCATAAATATACAGCCAATTATCGTTACAC tpg|BK006947.3|:730484-732411 7X163= 392=7X 
 tpg|BK006936.2| 328323 + tpg|BK006936.2| 328495 - INS TTGCTCATAGAATTCATCTTTGTCTTTAGAATTGACCTCATTTCAGTAGTCGAATAACCACTTTGAGTCTCATCTTTGTTTAACTTTTTAGATTTTTTGTAGATTAAAAGACGTGAGTTTTCATCAAACCTAACACTTGAGGTACTCCGATCCTTTATACAAAGATCTGTATCCATTTCTGAAATGTTTTCGCTGTCAGATAACTCTGCATCTTCTTCGTTATCAACATATGGATTGAAAGCATCATAGAATCTTTTATTTCTAAAATTCACGCATCTTTTCTTTTTTTGATGACTTTTGATCAAATGCGTTAAGTTATCTTGGCTTAAATCAGCTTTACCAACTTTTGAAAGAATTTGTGATATATTGGTCCTATTAGTAAGGCCGCGAAATGTGGGGATAGTATAAATTTTACTACTTCCACTTGAGCTTGTATCAGATAAATCGGAAAGTTCCTCAGATTCAACTGGCTCGAATGTGGTCTCTACATCATCCGAATAGCTACTGCTCGCATCATCTATGTCTTTATCCAATGTATCATCTTTTAAGGCCGAGCTCACTTCAATTGGTTTTTCCATTGCGTCCACCGTGCTAGTATTAGAGTCTGGTA tpg|BK006936.2|:327089-329729 7X440= 591=7X 
 tpg|BK006936.2| 741969 + tpg|BK006936.2| 742171 - INS GTGTAAAGAGTACCACATATATATATTGGATAGGATACTCTTCCGTTAAACGAATAATCGCCGTGTCTCAACGGGTCCTGCTTGGGACCCCCAACTTCACCAGTCTTGGGGTTAACATCACCTTCGAATTCAGGTATGGTCTTGGAAAATTCAGGCGAGAATGACCCAATATCGTTTTTGGTTAAAAGCGGTGAATTCAAACTCTCCTTTGTACGATCGCCGGTGGCCTGCGCATTATACTGATCTATTGCCTCTTGCGATGTGGCAATCCTCTGAAGTCTTTCGAACTCTTCCTGCTCTTCTCTTGGCAGCTTGGGAGGGCCGGGGATCCTTTCAGTAGTTATTTTTCGGGTGGCCATATTAAATGGTCGTCCACGGAGTAGATTTAAGGCTCCCGTGCGAGGATACCGATAACCTGTGCTTTTGATGGCGCACAACATTAGTT tpg|BK006936.2|:741065-743075 7X6=152S 12S342=1X67=7X 
 tpg|BK006947.3| 626640 + tpg|BK006947.3| 626908 - INS TTTCAGCTAATATAGACACGTATAGACACTCTTTTAATTCTTTCCTTTTCCCTAGAGGTAGCCAAAGTCTTTGCAACTATACTTTCAGCTCTGACAAATTTGTTCTTATTACTTCTCTTTTTTTTGATTTGTTCTTCCCTCTTTTTCTTAGCTAATTCTTGTCTTTCGATTCTAGTTCTATCAGCATTTCTTCTTTTCCTCAAAAGAATTTCTGGATTAGAATTAAGAGTTTGCGCTTTACTGTCTTGAGTTGAAGACATTGTGACTTGTATATCTTATTCTTTTTCCC tpg|BK006947.3|:626048-627500 7X3=262S 2S269=7X 
 tpg|BK006947.3| 714419 + tpg|BK006947.3| 714087 - INS AAAGGATTCTTTCCTTTAGTTCTTTCATGATTGGATCATTAATCTCTGGTGAGTATGGCGCTAGTAAGCCTGGTCCCTTGATTGTACCATCTAAGACGAATTTCGTTGCAATGGCAACTGGATAACCAACAGTAGCGGCCATAGAACTGTAACCACCAACCTTACCATAGTCAACTAAAGTGGATGTTCTTGTTTCGGTAGTTCCATCAGCCCATTCAATACCGAATTTGTGTTGTAGTACAACCATATCTCTTTCATTGTCTTCATATTGCATTAGTTCTTCTAAACGTGCACATAGAGTGTCTAAAGCATTACCTCTTGGTGTGATCTTTGCGTCAGAGAACAAGCCTAACCAAGCAAACCCGGAAAGGATTCTTTCTCTATCTTCATCATCTTTCCAAGTAGCCTTTGAGTCAATGGAAGCAATCAAATCTTCTTTAGAAGTAGACTTGGCACCTAAATATTGTTTTAGTGCTTCGTTC tpg|BK006947.3|:713109-715397 7X4=259S 467=7X 
 tpg|BK006947.3| 178451 + tpg|BK006947.3| 178526 - INS CTCATCAACAAATATAGACTTAGAACTTCAGCACATTGAATCTGAGATAAGTAGATTAGACGTTCAAAATGCAGAAGCTGAAAGGGACAAATATCAAGAGGAATCACTAAGACTAAGAACAAGATTTGAAAAGCTGAGCTCTGAAAACGCAGGTAAATTAGGTGAAATGAAACAATTACAGAATCAAATAGATTCATTGACTCATCAACTG tpg|BK006947.3|:178015-178962 150S60= 10S188=7X 
 tpg|BK006936.2| 578702 + tpg|BK006936.2| 578670 - INS GAGTACTGTCCTATTATTTGCCACTCTTCGTTCTGTATGTTACGAGGGCGTTCCTTAAAATGGGTAGACGCATCTTATTACCCGCCAAAAAACGTCAAAAGTTTTAGGAACACGTCTAAAAGTTGAAATAATATGTGAAAAAATTGATGAAATATTAATGAAATGGCTTATTTAAACGAATTCAAGTACAGGAAAGAGGTACGCACAACTACTTGAGTTTGCCAATATGTCCGAATTTAATGAAACAAAATTCTCCAACAAC tpg|BK006936.2|:578132-579240 7X3=349S 131=7X 
 tpg|BK006947.3| 223561 + tpg|BK006947.3| 223871 - INS TTCTTTATTCAATAACTTTTTTTTGATACCCCAGTATCACATTTTCTAACATTCGAAAATCCTCTTTCGATAAGGAGTTTTGTAGAAAAATTTTGGCACCGTTACAGTCTTCTAGCGAGATATCTGGCGATGTATGTTCATCAGTTGGTTGAGCAGAAGCCTGTTCATTTGCCCTCGTAAAATGCTTCGAAGAGTTTTCTCTAGGAGTAGAGTGTATGAAATTGGGTACATCCTTTTTATGAACATCAGTACCTATGGGAGACTTATCTTTTTCGTTTTTTGGTCGTTCTTGTAATCCTGGAGATTCCTGATAACTAGTATTTCTAGCATAATTCATTTGATCCATAGATGGTGATTTGTTCTCTTCATA tpg|BK006947.3|:222807-224625 7X96=1X471= 185=7X 
 tpg|BK006936.2| 476230 + tpg|BK006936.2| 476213 - INS TTCATTGTGTTCCTTGAGCTACCCTTTAAAGCTGGGGAGATGAGCTTGCCCTTCCTGTCATCGCCATTATGACGAGAAAAGTAAAACATGTAGAATAAGGTCCACCCAAACATGTCCGAGCAATGACGTTATATATCGTGTTCCCTGTTCAAAGCATGGCATATGTGCCATTAAAGGCGAATTTTTGTCCCTAGCAAAGGAGAGACAGCGAGCCACCATTAAGAAGTGACTTGAAAGCAAGCGAAAATAGCTACACATATA tpg|BK006936.2|:475677-476766 13S92=32S 126S5=7X 
 tpg|BK006947.3| 197852 + tpg|BK006947.3| 198626 - INS CTTATTCAACTACCATTGCTAGCTCCTCTCCGTGACGCTTATTCAGTGTCTGAACCAACTGCTTCCGCTTGAGACTGTTTTGCTCGCCATTGAGTAGGCCACCACCGTTCATGCATGCACCCGGACACGCGTTTACCTCGATGTAGTCCGAGTGGTAGGGATCGGCCGTGGCGGCCGTGGCGGCCGCCATCTCGCGTGAGTTCGCCTTTGGACCTGTTCGTCTCTTCCGCAGAGCGGTGATGTTCCTCTTGCGCTCTGACCCGGAGCCCGAGGTCAGTTTACGCACCAGATTTTGGATGTTTCTAAACCCGGAAAGCTCGCTGGCGGCGGCTATTATGCGATCATCGTGCAGCAATCGGTACTCGACAATGTCGCTGTTTCTACCCTCCAGAACTATCATCTGACTTCCTGGGTGTAGTCGTTGGACAGCCGTTACGTACTGG tpg|BK006947.3|:196952-199526 7X272= 430=7X 
 tpg|BK006936.2| 102649 + tpg|BK006936.2| 102771 - INS CTCTGCACTAAATGGCTACAAGACTCTGTAGGTGGTATGACGAAAACATGCAGTATCGCAACTATATCACCTGCGAAAATATCCATGGAAGAGACTGCAAGTACGCTAGAATATGCAACGAGAGCCAAATCAATTAAGAATACTCCACAAGTAAATCAGTCTTTATCGAAGGATACATGTCTCAAAGACTACATTCAAGAGATTGAAAAATTAAGAAATGATTTGAAAAATTCAAGAAACAAACAAGGTATATTTATAACTCAAGATCAGTTGGACCTTTACGAGAGCAATTCTATCTTGATT tpg|BK006936.2|:102029-103391 98S241= 9=1X24=1X250=7X 
 tpg|BK006936.2| 78077 + tpg|BK006936.2| 78325 - INS AATACCTCTAAACTATCACCTGAAAAATGCTACTGCTTTACTTGAACAAATTGTGGATGATCTTTCTATCGAGAAATTGAAAGAAGCTGTATCAATGATGCTGAGTGTAAATTATTACCCAAAATCTATTGAATTCTTATTGAATATTGCCAACTCTATGGACAAAGGCAAACTAGCTTGTCAATATGTGGCAAATGGATTTTTAGAAAATGATGATAGGAAACAATATTACGACAAACGTATCTTAGTTTATGACCTAGTTTTTGATACTTTAATAAAAGTAGACGAACTTGCCGAAAAAAAACAGTCATCAAAAACTCAAAACCAAATTTCGATATCGAATGACGATGAAGTGAAACTGAGACAAAAAAGTTATGAAGCCGCCCTAAAATATAACGATAGATTATTCCACTATCATATGTATGATTGGCTTGTGTCTCAGAACAGAGAGGAAAAACTATTAGATATTGAAACTCCATTCATACTC tpg|BK006936.2|:77089-79313 7X258= 244=7X 
 tpg|BK006947.3| 249580 + tpg|BK006947.3| 249504 - INS AAATAAAATAGTACGTAGTAATATTATTTAAATTGCATGCGTTTTTTTCGTTTTAAAAAGAGATTTTAGTGTGAAATGCAGTCAAAAGGTACTTTTGTCTGTTTTATAGTACTTGTACATCAGACAAGGATGAATTAATCTTTTTTAAAGCGGTCTCCTAGTCTCCTTCTGAAACCAAAAGTAGATCTCATTTCATCCCAAAATAAAAGCCTTAAAGCCTTAAATTTCTGTCGTGGAGTTGGCTTATAAAGATATTGAAAAGCAGTTGATTGGTCAGTGAAAGGATCTTCTTTAATAC tpg|BK006947.3|:248894-250190 12S168=1X96=9S 11S8=7X 
 tpg|BK006947.3| 267999 + tpg|BK006947.3| 268278 - INS AGAAGGGAGAAGACATTAAACCGTATGGAGGCAATGAATTTGAAGAGGTTAGGGAAGTGTTAATCGTGTTACCAATTTGCATCATTGGTTGTTGCGAGCTGGCAGAGAGTGCCTGGTTAGCACCATTATTGCTGGCTCCATTGTTGGAGCTGGCGTTTGCATTGGCACTGGTGTTGCTATTCGTAGGTGCAATGGCTGTCGATGCTGCAGAGGGT tpg|BK006947.3|:267555-268722 53S345=1X98= 108=7X 
 tpg|BK006947.3| 24033 + tpg|BK006947.3| 24607 - INS TGCTAGCTATACTTCCGTGTGACTTATTTCACAAAGAAGCTATCTACCTCGTCCATATCAAATACTGTCGAATTAACATATCCCGATGAAGGTACATCTGTCAGACTTTTAGGAAAGAGAGATACTTCAACCACCCTAGCCTCAGAATTATATTCTGAGTCAGCTGCTAACATTGATTCCACCACCAGTGATGACACAACTAGCTCTGATGCTGCTATAACACCAACATACTCAAATTCAACGCTTTCTTCTTATACTTCGCAATCATCCGCTATCCCTGAAGTTGCGGTTACTGCATCATTGAGTAGCGGGATCCTTTCTTCTACAGTTGACGGTGCTAGCACCTCGGCGGACGCTTCCATGTCCGCTGTCTCTACGGTTTCTTCTAGCAGTGAACAAGCTTCTTCTTCAAGTATTTCTTTATCGGCTCCAAGTTCTTCAAACTCAACCTTTACTACTCCTTCATCTTCTCTGTCTGCTACTGAAACATATAGTATTATCAGTTCAGCTAGTATATCTGTCACACAGGCTTCC tpg|BK006947.3|:22951-25689 7X364= 267=7X 
 tpg|BK006936.2| 141893 + tpg|BK006936.2| 141643 - INS AGTGTAGAGCCGGTGATAACATTCATTTGCCCCATATGTATTTTTTTTTTCTTTTGGTATAGCATTGATATATTGAAATTTGTATATATTGCTGCGAACACTATTTAAAACAGGTTTTTTTTTTATTTTGGCAGTTTGAAACCCTTTCCTCTGATGACTTTAGTGTAGTAAATGTAAAAGAAATCAGAGTACAACAGAGTTTGCAAAAGTCCCGCGAAGAAGGCAATCTTGTCCAATTTTTTATCTTCCGTGCTGTACCTCCAAATCCAGTTAGGAATATACAATGCTCTGTATAATCC tpg|BK006936.2|:141031-142505 7X191=1X115= 12S265=7X 
 tpg|BK006936.2| 136045 + tpg|BK006936.2| 136045 - INS CCCGAAGTATTTGAAGTATACTGCAAGCATCACCGAAACAGGAAATCACGAAGCTGACTCATCTGTGATTTTCCGTCCCCACCATAGTGATGTAACATGCAGTAACGCACGGCGGGCCGAAAGTCGGACTTTACCCCAGATTTGTAGTTGTATCCTATTGGATCACGGGCGACGGACAAGACCCGAAGTGCGGACCGGCATGGTCAGCTTGCACGGAAGCTTTAAGGGTTTCCCTTGTTTCGGCATTAGAAGAGGCATTTCGCACGTTTTACCGGGTCAGAAACTTCGAGGAAGCTGTGACAATTGGAAAAAAAGGCAAAACTAAATGCAATGTATCCGGTTGCCCATGCATTATTTGTGATGTTTTCGGATGTAGTTCGCTGCGCTCCGCGGCGATATATCCTCTAGCGAGAGGCATATGTATAAATATATATATATATATCTAACAAAAGCATTCAAGTTTCTTTCTCTGGTGTTACGTCTTTGTTCGACTTTCTCTGCTTACAGCCCTGTATGACC tpg|BK006936.2|:134993-137097 7X193= 260=7X 
 tpg|BK006936.2| 294140 + tpg|BK006936.2| 294470 - INS TCTTTCATTCCCTCGCTCAGATAAAATGGAATTTTGGGGCCTTGCTTGTTTTGTTGAATCTTATTAATGATCACCTTATGATTGCTACCAGTATATGGAGGCTTACCTACTAACATGTCATACAACAGACATCCCAAAGAATACCAATCACAATTCTGACTGTAAGCTTTACCTAATAATATTTCAGGCGCACAGTATTCAGG tpg|BK006936.2|:293720-294890 7X66=35S 8S1=159S 
 tpg|BK006947.3| 279215 + tpg|BK006947.3| 279172 - INS GATCTCTCGTGATTATCTTTTGGGTCATCACAAATTTCATCATCGTTGCTGTTGTCTTAGAAACCGGTGGGATTGCAGATTATATTGCTATGAAATCCATATCAACTGATGACACTTTAGAAACTGCAAAGAAGGCGGAAATTCCCTTAATGACCAGTAAGGCCTCAATTTATTTTAATGTAATTTTATGGTTAGTTGCATTATCGGCATTAATAAGGTTCATTGG tpg|BK006947.3|:278706-279681 7X62=51S 2S1=233S 
 tpg|BK006947.3| 158333 + tpg|BK006947.3| 158967 - INS CCTATCCTACGAAGCATCATCTATATTTTCGTCAATTGCCCAGGCTTCATCCCAGGCATTTTCTTCTTCTTCTGGTTCTTTTTCCTTCTCTTGATTTGTTTTTTCTTCCTCGTCGTCAATATTTACATCAATTTCATCACCCCATGCATCGGCATCATCATCCTCTACTTCCCAATTCCAATCATCATCTTTGGATACGGCATTATGGAGTTCTTTTTCGTTCTGTACATCTGAATCATTTTTTCCAATTTTTTCGCTCATCGTATTAGTATTGCTAGTAGTGAGCTCAACTACTTCCAAATTTTGCCAGCTCTTTTTTGGATCTTCAAATATACTTCTTATCTCACTAATATGCGATTCAAGAACTTTATCTAGTAATAAATTGTAGTATAATTG tpg|BK006947.3|:157527-159773 7X190= 372=7X 
 tpg|BK006947.3| 194039 + tpg|BK006947.3| 193940 - INS TGTCTGGACTGCATTTGGTAGACAGTTTTCTCGACAAAACTCACGAGTTCAACAATGGTGCCAGAAGTAAACTATCCTCTCAAGGTTCATATGAAATGGACAGTTCCTCTGGAACTGCCACAGGTGGTATTTTACTTCCCCATGAGAGTTATCTAGACTCTGCTCAGCCAAAAGAAGAAGATACTCCACCAATCGCCTCAAAAGAGCAAGAAAGGGATGTGGATATAAGGGGTAGTATAGATG tpg|BK006947.3|:193440-194539 7X207= 228=7X 
 tpg|BK006947.3| 142002 + tpg|BK006947.3| 142730 - INS TATCAGAAAGTACCAAACAAATCCGCGCTCAAATTATTTCATCAATGAAGGAGGTGCAGGATAAATTTGGTTACCATGATTTGGAAGCCCTTCATGGAATGGCAGGTGAGAGAAAATTGGAAAACGATTTAATGACGGGTGGTATTGACACTTCATATCTAGGTGAAGATTGGGCTACCAAGAAAGAGAGGATACGT tpg|BK006947.3|:141594-143138 7X127=20S 1S1=164S 
 tpg|BK006936.2| 626202 + tpg|BK006936.2| 626903 - INS GGCAGGGCACACAGTTTGTCCGTCAACACAAGAAGAAATTTGCGTCTTTCAGTCTGACTTCTGATGTAGAAGAGAGAGTTATGGAATTAATCACCTCTGGTGATGTTTATAATAGGCTGGCAAAATCTATTGCACCGGAAATCTACGGTAACTTGGACGTAAAGAAAGCGTTGCTGCTATTACTTGTCGGAGGTGTTGATAAAAGGGTAGGTGACGGTATGAAAATCAGAGGTGATATCAATGTTTGTCTGATGGGTGATCCCGGTGTTGCCAAATCTCAACTGCTGAAGGCCATTTGCAAAATATCACCTCGAGGAGTGTATACCACTGGTAAGGGTTCCTCAGGCGTTGGTCTGACCGCTGCCGTCATGAAAGATCCTGTCACGGATGAAATGATTCTAGAAGGTGGTGCCTTAGTACTCGCTGATAACGGTATTTGTTGTATCGATGAATTTGATAAGATGGATGAAAGTGACAGAACGGCAATCCATGAAGTTATGGAACAACAAACAATTTCGATATCCAAGGCGGGTATCAATACAACTTTGAACGCCAGAACCTCAATCTTAGCGGCAGCAAATCCGTTGTATGGTAGATATAATCCTAGATTATCACCTCTGGACAATATAAATCTACCAGCTGCTTTACTATCCAGATTTGATATTCTCTTCTTAATGTTAGATATACCAAGTAG tpg|BK006936.2|:624800-628305 7X211= 684=7X 
 tpg|BK006947.3| 770849 + tpg|BK006947.3| 771081 - INS GAATAACCTTGCTTGGTGTGTGCGATCATCCAACAATTTAAATTCAACAACGTAAACGCCCTTGTAAGGATTCTCAACAGGGGACGCCTTGTACTGCTTAAGATTTAAGGAACTGATACTGCTGTGATTTGTGTTACCACAATTGTTAACAGTTAACTTGTGAGGACCATCATCCAGGCTGAAAACACCCTTGGCGATACGGTTGGCATAACGACCAACTGTAGCGCCCATCATGTTACCATCTGTTAAATAGTCTTGTACGTTTGAATAACCTTGAACGACTGATTGGCCGTTTACCTTCAGGTCTACCAAAGTTGCACCAAGTGGCGCAATGGTAGCTTGGAACTTTTTCTCATCACCAATTGTAATG tpg|BK006947.3|:770095-771835 7X224= 41=1X305=7X 
 tpg|BK006936.2| 523009 + tpg|BK006936.2| 522478 - INS AATGATAAGCTGTGCTCTTGTTAATAGATTTGGATTATTCAACCATTGACATTGTTTTGAAATAAAGAAATTCATTTTTTTCGTTAACTCGAGTTTAAGACTTTTGTGCACCTCATAAGCGGGATTTCGTGACTCAAATGATAAGCTGTCTCCTTCATTATCTGGAGCGCTCTTGCTTTTTTCCAACTCTTGCATATCAGACAGAATACCTGACATAGAAGCTAGAATGCCTGCCAAGCTTCTAAAATCTACTAGTTCCTCTTGCGTAACTGATTTCGAACAGCTGAAGTAAAACCACTTCTTGTAAATCACGTCCATTGAATCCAAAAGGATTGAGTCGGATCCTTTGATATAAGTTAAAATATTATTTCTTAGACGCCGTGGCAAAGCCACTGATCCTGAGGCAGTGAAATTGTCCTGGGCCATAGCATCTATGAAATCAATATTGTAAATGGAATATTGATCCAAAGCGCCTACGTATTTTTGATAAAATCTCAAGGATCGTAGAAATTCACAACATGAAATTTTTATTAAGCGTGGCGTATTTCCACGACTGCAGTATAATGAAATGAAAATTCCACTTCCTACAGCACCAACTAATAATGGCAGCGTCAACCTCTCCGTCGTAATTATTGCCTGGACTAGGT tpg|BK006936.2|:521170-524317 7X5=393S 362=1X264=7X 
 tpg|BK006936.2| 778784 + tpg|BK006936.2| 778879 - INS CCCTTGAAGTTCTTATAGACCTCTAAAAAGGTAAAACAATCAAGCGGGCCTTTTGACTTCGAAGTGGAGGCTAAGCACCAATAATTGAGCTTATTTATAACTGAGAAATACTTATAGACCTCTAAATCTCTTCCAACCATTGAATGGTCTAAATAATCATCACTACTGCTATCTTCGAGCAATTGAGGACATGTGGACTGAACGCGGGTCCACAGGTGCTTGAAGGAGGGAGCTGTTGCAC tpg|BK006936.2|:778288-779375 27S100= 94=34S 
 tpg|BK006936.2| 667478 + tpg|BK006936.2| 667722 - INS TTGGTACTTAACAAAGGCACCGTTTTTGGAGTGGAGGTGGGACCACTGGTATGCAAAATCAGGGCAACGTCACTGGAACGGGCAAACCCAGGGAATTTAACGGGATTTGTGTTGACAAATTTGGCGTTGTTCAAAGACCGGTAAATAACCCTTTTGTAGTTGTCCTCTGGAGAGTATATATCATACTCTACCCTAAACCTGGTCGCATCGAAGGCCAGCTCTACGATAAAACATCCAAACGTGGAGGCAGATTTTAGAATTTCAGAACTCTGTAACTTTGTGGTACCCTTTGGGACGCAAATCGCCTTAGATTTCAGGTCATTCAAATAAAAATTGAACTCCTTTTCCTTAGAATTGGGATTCAAGGGCGCGCCAATTTTAGCGTCCATAGTAACACCGAGGAAAGCGACGATAAATTCCAGCCCATTACGCATGGATATCGCCACTGTATCTTGTCTGAAAACAGCTCCGTACAATGGAGAATTAGGATTTGTGAACATGGTCTGGAAGTGACCCACCATGTGGGATAGATCCCTGTAGGTC tpg|BK006936.2|:666378-668822 7X305=4S 24=1X310=1X41=1X149=7X 
 tpg|BK006936.2| 560834 + tpg|BK006936.2| 561491 - INS TTCTATGAGTGCGAAGCGGATGCAATACGGTATTTCATCCTTTCGCATTATGGTGGTATTTACATTGACTTGGATGATGGTTGTGAAAGAAGGCTAGACCCTTTGTTGAAAGTACCAGCATTTCTAAGGAAAACTTCGCCTACAGGAGTGTCAAATGATGTGATGGGCTCTGTTCCAAGG tpg|BK006936.2|:560460-561865 7X10=80S 85S5=7X 
 tpg|BK006947.3| 355079 + tpg|BK006947.3| 355373 - INS AAAATAAAAAATGGGCCTCGGCGGAATTTGAATTCGGGTTACGTTTCCCACGGAGCCCCGGATAGAAAAGATTAGTTTCAGGTACATGTGTCAAATGAGGATAAATCTCAAACACCCATGTACCGAAAATCGATGTGTTGGTTATATTACAAGGTTGGAATAGACCACGGTGATAAGACGTGGAATTTTTGACTGACCATGCGACTCTGAAGGTGTTAACCGG tpg|BK006947.3|:354619-355833 7X11=1X174=16S 2S1=210S 
 tpg|BK006947.3| 259033 + tpg|BK006947.3| 259279 - INS GTTTTTACTTTTATAAGAGGTATAAGAGTAAGGCTCCAAATCAAAGAAAATCTAAATTTGAAAAGAAGTTCGTAATTTCTAATATTTACACTTTTAGAGTTTGGGAGGTCGTATGTTCGAGTCATGGATACTATGAATACAGCAAACACTTTGGACGGCAAATTCGTTACTGAGGGTTCTTGGAGACCTGATTTATTTAAGGGTAAAGTGGCATTTGTCACTGGTGGAGCTGGCACGATATGTCGGGTACAGAC tpg|BK006947.3|:258511-259801 15S183=11S 2S237=7X 
 tpg|BK006936.2| 595913 + tpg|BK006936.2| 596673 - INS AGTGCATTCCGAAGTATCCACTTGCCAAAAGAAATCTCAAGGCTTCAATGGCGCTCGGCGCAATTTTGTTCTTATCTGGCTACATTTCGTGGCTACTTGATATACACTATTGTTCGTTCTGGGTGCACGTTAGAAGAAGTATTTTGGCTTTACCACTTGGTGTACTGCTTGAACC tpg|BK006936.2|:595549-597037 192S20= 154=7X 
 tpg|BK006947.3| 117668 + tpg|BK006947.3| 118285 - INS AAAATTGAATCTCCCGAAGGCCACAATGCCTTCCTATTGGAGTTTAAGCTGATAAACAAACTGATAGTACAATTTTTAAAAACCAACTGCAAGGCCATTACCGATGCCGCTCCAAGAGCGTGGGGAGGTGACGTTGGTAACGATGAAACGAAGACGTCTGTCTTTGGTGAGGCCGAAGAAGTTACCAACTGGTAGGGATAGATACCACAC tpg|BK006947.3|:117234-118719 7X24=1X80=52S 5S1=331S 
 tpg|BK006936.2| 576009 + tpg|BK006936.2| 576194 - INS TCTTACAGTCTCCTCGTATGATGTGATTTTTGGTAAGGGGACGTTCCAGAAACGTCTACTATTTTGGATGATTTACATAGTTTTAAAATAAAAAAGGCTCAATTTTACCTTCCGCGCATTTCTATTTTTTTAATCTAAAACCTCAAATCTTACAGTCTCTCCTAGCCGCTTTCCTGAAGGATCATGACTAACGTTTGCCAACCAGCCGATGAGACAAGTTTTAGTAGAGATTCTTCCCATTCATTTTTCACAGCAGATTCTATTAGTA tpg|BK006936.2|:575459-576744 7X279= 30=1X221=7X 
 tpg|BK006936.2| 734026 + tpg|BK006936.2| 734531 - INS TGCCACCATCTGACCTTGTGACCGAAGAATCCGTTTCGTCGAAATCATCGGTATCTGTAGGTGTGTTATTTTCTTTGACCACGATTGTCCCATTAGGTTGCAAACCAACAATACATCTTTTCAGGAATGCGACGAGTTCTGCATCTGGCAGGTGTCCCACGCACCATTGGCACCAGATCAGCCAGTACTTGCCGGCATCGGGGGTCCAGTCCTGCATCCCTACTTCATATATTTGTCCAATTTGGCCTTTGTCTTTCAGCTCAGCCAATTCAACGTGCATTTGCTCGATAAAAGGCTTTACCGGTTCTACAA tpg|BK006936.2|:733388-735169 13S216=51S 34S5=7X 
 tpg|BK006947.3| 545655 + tpg|BK006947.3| 545852 - INS GGCTTTGAACACTGAGTTTGGAACTATCAGCCGTCAAATACGCATAAAATAACATCAAATACTCCAATAATGAATCAGTTAGGAGCTTTAGCCGTAAGTTCTAAATTGTAAACACATTTGCATCATTGAAAAACTATACTAACGCGTTAAC tpg|BK006947.3|:545339-546168 7X1=2I10=62S 66S10=7X 
 tpg|BK006936.2| 648240 + tpg|BK006936.2| 648039 - INS TTCGTTCTCCCACTCAAAAGGATCATCTACTTTACAAAGTTCTATACCATCTACCCCAGAATTTTCCTTGTTTGTTGGTGATCTTTCTCCCACCGCCACTGAAGCTGATTTGTTATCTCTTTTCCAAACGAGGTTCAAATCTGTTAAAACCGTCCGCGTGATGACTGACCCTTTAACAGGATCATCTCGTTGTTTTGGATTTGTCAGATTCGGTGATGAAGATGAGCGCCGCAGGGCACTGATTGAGATGAGTGGGAAATGGTTTCAAGGAAGGGCCTTAAG tpg|BK006936.2|:647461-648818 7X345= 9S256=7X 
 tpg|BK006936.2| 501986 + tpg|BK006936.2| 502200 - INS GTTACCGCCACAGACATATTTTCTTCTCGTCTGGTATTCATCAACGTTTCTTCGCTAAATTTTAAACGGACTGTGCTGTCATTGGGCAAAGTTGACAAGAATATATTGTTATATAAGTTTGCCGAGAAGAATCCGATAAAGCCATGGATTTCGCCGCGGTGCTTTATCTTGAACTCATTTAATGAACTTTGAGAAAATTCAACTGTAAAATCATCTTCGTCTTGGACAGTATCTTTTTGGGCCATGGGATGCTCGAACCGCCACACTTCATTTACCCTTGAGGATAATATACAGTATGGCACTCTATGGACTATCCAGGGCGCCTCCAAAGAGCGATTTGTTTGTGAGAGTTTTTGGTAGAATAATGGTGACGAAATGGGTGCTATGTATGAAGAGTATGACCTCGGTATGAAAATTGTGTCATTGTGGGAATGATATTTTTCAATAGACCAGAGACATTCTGGTGATAATTCATTGCAACCGAACGAACCCAGCAGTTCACTTATGCACAGATCTATCT tpg|BK006936.2|:500932-503254 7X255= 1S503=7X 
 tpg|BK006936.2| 503428 + tpg|BK006936.2| 503843 - INS GCTACTAGGAGGCGCCAATATTAGCTTATTGATTCCAACAAACCTCGCGTACTTACATTCGTTTAGAAGGACCTTTAAGCCAAGATCTCTTACATTTGGATCGCGACTCTCCAGCTCCAGCCAAGAGGATAACAGCCCTATGTAAGACGGCGTATCGTCATTGTCTAGCTTCTTGACGTTGAACGGGGGTATACAG tpg|BK006936.2|:503022-504249 7X6=289S 98=7X 
 tpg|BK006947.3| 447516 + tpg|BK006947.3| 447545 - INS TCGTGATCCTACTTGCCTATGGACATTGAAACTTGGCTATAAGTTCCGTCAAAGGGGGAAAAAATTGCTTTGGAGAAGGAATAAAAAGATGAATAGTCAAGGTTACGATGAAAGCTCTTCCTCTACTGCTGCTACTAGCGGTCCTACTTCTGGAGACCCACGAATGGGTAAGAAACAACGGTTTATGAATCTCATAAGAACCACAAAGGATGTTTATATTCCTAACCTGACGTCATCCATTTCTCAAAAGACAATGGATGGCATCAGGAGCACTAC tpg|BK006947.3|:446950-448111 77S291= 3S256=7X 
 tpg|BK006945.2| 684486 + tpg|BK006945.2| 685107 - INS GCCTTGGTTCCTTAGAAAACCCTTTTTCGGAGTCACGGTTGTTCACATTTTGTTCTTTCTGCATACTGGCCTTCGATGCAGAATTGTAAATAGCCCAAAGGATATTAATGACATGTTGATCAATCAATTTTTGTTCATACATCATTCCTAATAGCTGTTCCAAAGAGGCCAAGTCTGCAATAGATGCGCCGATGCTTAGATTAATTAAATTTTTGGCAATATGTGCCGCCTTCTCCTGCATATTGCAACTATCTGGCGCGGTTAAAAATAGCTGCTTATAACATTCTATCAAATGTACTGATATACTCGTTCCTTCATCGTTTGTGCCCTTCATCCAAACCAAATGCAGCATTTTTTTTATACCAAATTCGCTTAACTCAATGTC tpg|BK006945.2|:683702-685891 7X161= 193=7X 
 tpg|BK006945.2| 828042 + tpg|BK006945.2| 828295 - INS CCCCGGCATTGAGCATCGCATGGATGAGTATGGCGTATTTTGATTGCTCATATATAGTGGGGGGGAATACTCATGCTGTGAAAAGCACAACTCTTTTCACTCAACGAGGTTAATGCCTTCTTTGTCTCCACGCCGTTTTTTTCTGGCGCCCTTTTGAGAAAGATAGCCTGTCCCGTAATCGTGGCTTTGGCAGAGACAGAGGGTGAGCGAAAGAGCGGGCGAAACCGAGAATGGATTCCGAGTAAAGGATTGCGATGGCATGAAACAAAACCGAGAGGCACTCCTTGTAAGGACACACATACACAGACGTAAACATATATATACATACGTATACTCAAATATATCTTCGTATCATTAGGTCAGCTTCTCTCTTCCGCACGTAGAATTAGAGAATTAACGCAAGACTATACCATTATAAAAACGCATAAGAAACAGTTTCATCATGATTGACCGCACTAAAAACGAATCTCCAGCTTTTGAAGAGTCTCCGCT tpg|BK006945.2|:827044-829293 7X243= 477=7X 
 tpg|BK006936.2| 234630 + tpg|BK006936.2| 234090 - INS TCGGTATCCAAATTATAATGATAATGCATCCTTTTTAAATCTTGGGTTGAGAACTTATAAGGTCTACTTGAAAAGTATTGGGTTTGAACATACTATTGAGCTAGACGAGCTTGCCATCAAGCGTATAAGGTACATTTTGAGCGATACGTCGGTAGGATCAGAACATCAGTGGGATTTGGTATACTCAGCTTTAAATACGTTCTCATCTTATATGGAAGCAACAGAGAGCGTTTATAAACATGGTTTCAAAGACATATGGGATGGTATTATCACATGTCTCTTGTATCCGCACTCATGGGTCCGTCAATCGGCGGCAAATCTTGTTCATCAACTCATAGCCAATAAGGATAAGCTGGAGATATCATTAACCAATCTGGAAATTCAAACCATTGCAACAAGAATTCTTCACCAATTAGGTGCGCCTTCTATTCCGGAGAATCTTGCGAACGTCTCAATAAAAACATTAGTTAATATCAGTATCCTATGGAAGGAGCAACGCACGCCGTTCATAAT tpg|BK006936.2|:233050-235670 7X205=12S 2S495=7X 
 tpg|BK006947.3| 324631 + tpg|BK006947.3| 324350 - INS GTGTCATAGACTCCCAATGCGATAAACCTCCATTAAACTCATAAGTGGTCTCTCGAATAAACGAAAATGTCTCCATATATAAATATGAATTCTGCACTATTCTAAAAAAAATGGAAAGCCATAATTTTTCGAGCAGGGTAGAGCACGATTTTATATTTCATAGAAAAGATGAACCTGATGTTCATATCCCCATGATTAATTACAATCAAAGGAAAAATGCGGATACGGCAATTCATGGATTAAATCTTCGTTGGTACGGGACAACTAGTTTAGCTTCACCTTTTGGCTCAAATAGCATCAACCTACTTGTACTCGATGATACGATGGCATCCTACATGAACCAACAAACTATTGAAGAGTTTGATTCTTACAGCCGTTCCCGTCCCACAAGACCGCTGGGTTATCTCCCAGTATGGGCCAGATACACAGA tpg|BK006947.3|:323476-325505 7X165= 215=7X 
 tpg|BK006936.2| 551725 + tpg|BK006936.2| 552083 - INS GAGAAATTATTTTTGGTTATTTTATTTCTTACTGAGAATATATCTCTTAACGCTTCTTGCATATCAGTATCCGTGGAGTTTATTGACTTAAACTTTTGAGAAACTTTTTTCATGGGGGAGCCTGTTAAATCGATTGATGAAGAGGAGTATTTGTGACCAACGTTTCCACGGGAAATTTTGTTTTCAAATGATTTTGTTGGAATAGATGATAGCCTATCGAAAACACTGGATGCTTTTGTAGATCCCGCGGTATCACTGTTTTCCACAGCTCTTATAGCAGGACTATTTATCGTAGATTTTTTTTTAAATGCGATTGGTGATTCCTTTACTG tpg|BK006936.2|:551049-552759 7X164= 166=7X 
 tpg|BK006936.2| 383984 + tpg|BK006936.2| 384098 - INS ATGTACAGGAAGCCTACTACCAAAAAGCACAAGACTTGGAGTGGTGATGGCTACGCTACCTTAAAAGCCAGTAGCGATAAGTTATGCTTTTATAACGAAGCAGGGAAATTTCTTGGGTCAAGTATGCTACCAAGTGATTC tpg|BK006936.2|:383690-384392 7X5=65S 65S5=7X 
 tpg|BK006945.2| 223446 + tpg|BK006945.2| 224188 - INS CCTTGACAAATACTATATTATTATCTTTTAGTAGGTCCCAGGAAGTGCCTTATTCTCAACATGTTCAGCGTTTATCTTTCTCAGCCTGAATGTATTTCAAACGATGACTAGAAGAGATTAGTACCCCTTATATAATCCTCGAAAATGTTGCTATCTCAGTGAATTGAAAGTTCATGCTGACGTCTTTATCAGCGTTATCCATTGCCTTGTTCTTTTCAGTGCAGTGGCAGATGTTACGAGGG tpg|BK006945.2|:222948-224686 243S294= 121=7X 
 tpg|BK006936.2| 651652 + tpg|BK006936.2| 650933 - INS AGCAACACATACCGCTGGAGGACGCTGTCGTCAAACTAGGTGAGCTGAGAAGAGGAATTAGGCTGCTGGCACCAGACGACAAGGATGTCAAGTACCGCATGGATTGGGCCAGACGCTGCACAGACCTCTTCGGCATTCAGCACTGCCACAACATCGACGTAAAACGTCTGCTGGATCTTTTCAAGGTCATGTTTCAAGAACAGAACTGTTCCTTGCAGTTCCCTCCCAGAGAACGGTTGCTTAGCGAGTACTGCTCGTCTTGAGCAACAGGGCCTCCTCTTTTAAGG tpg|BK006936.2|:650345-652240 7X5=183S 248=1X21=7X 
 tpg|BK006947.3| 484278 + tpg|BK006947.3| 484139 - INS AAGCAGATCAGTACTATAGAAGACAATGGGACAAGCTTTTATTTGCCAAAAATCAACAGAATCTTGACTCAACGAAATCATCTGTTTCATCAGCGAACACAATCAACTCAAACACATCCCATGATCCCGTACGAAAAAGTTTACTCAGTGGACTAT tpg|BK006947.3|:483813-484604 7X82=35S 1S1=173S 
 tpg|BK006945.2| 260044 + tpg|BK006945.2| 260038 - INS TTTGAACAAGCGGTCCATATGTACACTATTGCCTGCCAAGACGCCAACGTTCTTGTCTGGGATGTAGCGCTGGATGTACTCGAGCAGCTCATCTTCTACCTGGGCCAAAGTCTTCTCACTTGCCAAAACTTTGGCGGTGAGACCGCTATTACCGTGGTGCTCAATACACCACTCGTTCATTTTGTTCATCACCTCGGGACCATAATGGATGACGCTCTCATAATGCGAGTCTCCTTGGCCATCGGCCGCTTTGACGGGTGCCAGGTGTCCATCGGTGATGATGCAGCAAATCTCGATAATTCTGTCATTCACGTGGTCTAAACCGGTCATCTCGCAGTCGATCCAGACCAAGGGTTTGAACAGCTTGGTTTTAAGTTCGGGTGTTTGCGCCATTGATTGCAGGTTTTGGATGGTTCGAGGACGTAAGTACTGTGAAACGGATCTTCTGTACAGCGAGAAGAGGTTTGGG tpg|BK006945.2|:259086-260996 7X8=143S 235=7X 
 tpg|BK006947.3| 221938 + tpg|BK006947.3| 221636 - INS CTGGGTTCTTCTGCACCTTCTTTCATTCTTTTATCGAGCTTTTTTATGAAAACTACAAACCTTTTCACGGTTTTGTTGTATTCATTTCGAGCTTGTTGCCTAGCCTTCTCATTTCTTCTATTAACTTCCCTCTTGGTTCTTCTGTCATAGTTTTTAGAGTACATGTACTCGTCTTTCCAGCTAAAACTTTTCAAGGTATTGAACGCTGACCAAGTCTTATAGAAATGTTTCAAATATTCATAATCCGTTGGCGAATATCCAAATAAAGGATATAAAAGTTTATCCGTCTTGTTAATAAAGTTATCGCAGGCTTTCAAATAGCCAATACTATTAATATCCTGTTCGAATACATCATCTTGATACTCGGAAAATTTCCCCAGTCGCTTACCACTTAAAATCTCATCTTTAGCTAACTTGGCAAATATTTTTCCTGCAATTTGATATATCCCAGCAGCTGAGTTGTCTATTTTAGTATAAAGAGCAGAGTTAAAAAATAAGAGTAATTCATCAGTTGTGACACCTGTGACTGTAGCGTCTACCTCATAATCATAGTAATCATCAGTGCTTGGTGGAGTATCATTTAAAATTTGTTCCTTATGTGAGTCATACCATGCTCTTTCCTGGGGGTCAGACAGTACTTCATAAGCGGCTCGAATCACAGCAAATTTTTGTGTGGCTTCTTCAACATTATCT tpg|BK006947.3|:220236-223338 7X14= 672=7X 
 tpg|BK006936.2| 43445 + tpg|BK006936.2| 44115 - INS GTCAAAGAGATTATTCCGTGTTAATTAATATTCTATATTCAAAAAAGTTAAACATATATACTGCATGTACTTACCGCCGAAGCACAAACGTGCCACTTCCATGAACACTTGCTCTTTATTTATAGTGGGGCTGATATGCGATGGCGTAAAGCTACTCCAGCCTCCTTCTTGTCATATCCTCATGACTGTCACTATGTGTTGGTGTAGCCATCGAACTTCCACTAGATTTGTTCTTCCTTTTCTTACTATTGTTACCTGAATTTGAGCCGGATTGGCTTTTTCCTGTACCGTCTAGATC tpg|BK006936.2|:42835-44725 7X5=193S 152=1X127=7X 
 tpg|BK006936.2| 22524 + tpg|BK006936.2| 22634 - INS AAGTGTGTCTATGCTACCATGCCTAAAAGAAGATGAAAGGAAACTTCCTGCACGAAATGACGATGATGGTGATCTTACCTTTGGGGAATATGTGGAAGATACGGATGCTGGGCCCAAGCTTTGTGGATTATAAGAAAATGATGATGAATATGTGTTTGGTGTCATCATATCAGAATTGATGCTAGAAGATAAAGAGGAGCTCAAATCATCAGTTAAGTTATACATTGTGTCATCGGTGCCATGCTGAAATAAAAAGTCATGTGGTAACTCAGCTTTTAAGCCTTCTTGTTGCTGTAATGGAGTATTCATTGCTCTATCCACAGGTGAGTCGTAAGCCATAGAATAAGATGATCTCAAGGGACCCTGCCCTATGG tpg|BK006936.2|:21762-23396 7X13=1X119= 187=7X 
 tpg|BK006936.2| 285769 + tpg|BK006936.2| 285807 - INS CTTCACCATCAGAGGAAGTCGCTTTATTCCAAAACATCGAGGATGTAGGCAACAAAGTAGATGGATTACGGGAATGTACAGCTTTGTTTTCATTCGAGAGTTTCCAAGCATTTTGAGTGGTCATTGTTGTCATTCCTCTGTATGAACCAGAAGATTGTAGTGAACTGCTCATGGAGGTGTCTAGATCTATCACAGATTCGTTAAATTGAAACATTTTGGAGCTGTGTTTTTTCAGCAAGTCAAAGGTTGAAGCACGCTTGTGTCCCAACGACTTTTTTGAGTATTTCTTTGGCCTCAAATGAGGATCTACTTCCTTTAGAGG tpg|BK006936.2|:285111-286465 7X175= 302=7X 
 tpg|BK006945.2| 528660 + tpg|BK006945.2| 528966 - INS GTTTAAAGATCTATTCAGAACTTATGAAAGGTGCTGGTGCGGCTGCCAGGGTTTTTGAATTAAATGACCGTAAGCCATTGATTCGTCCGACTATTGGAAAGGATCCTGTGTCATTAGCCCAAAAACCCATCGTTTTCAAAAACGTGTCATTCACTTATCCCACTCGGCCCAAACACCAGATTTTCAAGGATTTGAATATTGCTATCAAGCCTGGTGAACACGTTTGCGC tpg|BK006945.2|:528188-529438 7X9=105S 109S6=7X 
 tpg|BK006936.2| 565905 + tpg|BK006936.2| 566119 - INS CAGCATTACATGCAGAAATAGCAGGGTGCAGAGGTCGAAGTAGATAGAGGACAACACCTGCGATGGCCGTACAGACACCAAGACAAAGACTGGCTAATGCCAAGTTTAACAAGAATAACGAAAAGTATAGAAAATACGGTAAGAAGAAGGAGGGCAAAACTGAGAAAACCGCACCTGTGATATCCAAAACTTGGTTGGGTATTCTTCTGTTTCTTCTCGTAGGTGGTGGTGTTTTGCAACTAATCAGCTATATCCTATGAAGCAGTGGCAAATTGCATATATAAGTGTACAGTGGAAGCAAGTACGTAAATAAATAAGCGATTTCGAATAATAATAACAACAAGCATAAGGCAGTATTACCCG tpg|BK006936.2|:565165-566859 7X3=266S 182=7X 
 tpg|BK006947.3| 122665 + tpg|BK006947.3| 123020 - INS CTCTCTATGGTGAGCTAAAGAAGCATCAATTGGTATACAAGAAAACGATTCTGTCTATGGAAAGTGGTAAAGTGTTAAGAGCTGCCATTAGATTGGCTCTGGATGTTATCAAAATCGACCGATTATCAAGAACTCCTAGGGACAATATGGTTCTCAAATTGGTTTTGAATTTTTTCAGAAATGTCATTGCTATAGAACCCGGTGAATTTACTATCAATACTAAGA tpg|BK006947.3|:122201-123484 7X151=17S 1S1=274S 
 tpg|BK006947.3| 765100 + tpg|BK006947.3| 765108 - INS TTAAATAAGCTTCTGAACAAGGGATTCATCTTCGTAAGGCAGGTGTAGCCATGGAATGCGTTTCAGTAGAAGGTTTGGATTCTTCTTTTTTGGAGGGCCAAACCTTTGGCGATATTTTGTGTTTACCATGGACAATTATCAAGGGTATCCGTGAGCGGAAGAATCGCAATAAGATGA tpg|BK006947.3|:764732-765476 7X152=13S 1=155S 
 tpg|BK006947.3| 607450 + tpg|BK006947.3| 607656 - INS GGCTGTTCTGAAGGACGCTGACATTCTACTATTGGATGAACCAACAAATCATCTAGACACTGTTAATGTGGAGTGGCTGGTAAATTATTTGAATACTTGCGGAATTACATCGGTGATTGTCTCTCATGATTCTGGTTTTCTGGATAAGGTTTGTCAATACATCATACATTATGAGGG tpg|BK006947.3|:607082-608024 7X39=49S 4S1=316S 
 tpg|BK006947.3| 347571 + tpg|BK006947.3| 347600 - INS GAGTATGACTATGTTCATGGTTCTACGATGAGACAGATTACTCCCCAGTGTGTTAGCACAAGTCACGAGGATAAGGATGAGGGACAGCCCTACAGAAATGGCAATGTTTTCTCCATGTCATCTAAATCAGATACAGCGGTATTGGCAAATAGTAATGACCCAATAATTTTACCTCCAACTTTTTCAGCATCCATGGGTACAACGTCTACATTAGAAA tpg|BK006947.3|:347123-348048 7X4=104S 104S5=7X 
 tpg|BK006936.2| 403335 + tpg|BK006936.2| 403450 - INS CCATGGACACCTTGCCATTCTCTTTGGCCAACATATGAGCTCCCATATTCAATCCTTTTCTTCCAGAACCAGCAACTTCCTCTTCCTCATCTAATTCGTAGTCTTTGTCTTTTTCCATATCTTCAATTTCCTTTTCTAAATCAGCCCTGTTTCGGATTGTGATATTTGGAATCATGCGAATCAACTGAAGAGATTTCTTCTGCATAGCAATAGCATGCCCTCTCAAAAAATGTGAAGGATCTGAATTATAGGTCAAACAATTTTTCCATATTAGCATAATATCGTCTACAAATTCTTGTTTGGAGTCATATTGAAAGC tpg|BK006936.2|:402685-404100 7X181= 159=7X 
 tpg|BK006947.3| 146239 + tpg|BK006947.3| 146589 - INS AAATTGAACTTGACGGATCTTAGTAGGAATACGCCAAAGGCAATAAATAAGTAAAATTTTATCAAAATATTCAGGTTAAATGGCATGGTCACGTTGGTCAAAAGCTGGGCGAGAATCAATGGAACAAATTTGTAGCCGACATAGCACAACAG tpg|BK006947.3|:145921-146907 7X7=69S 72S4=7X 
 tpg|BK006936.2| 729566 + tpg|BK006936.2| 729801 - INS CTCTTATATAGAAAAATAAGACAAAAAAAAAGGCCATCATATTTATACAACGAAAAGTGTTTAATATGGAAGCAGCAAGCGGTATATGAACTCAGTTTTAAGGTGTAGTTTATTTTATAGTCATGTCCATTGACGAGGCTGTTGCCAGATATAGAGATGTTATAGGCAATCTAGCAA tpg|BK006936.2|:729198-730169 7X5=83S 84S5=7X 
 tpg|BK006936.2| 719423 + tpg|BK006936.2| 718973 - INS GTCAGTTGAGAGTATTGCTATGATTCACTACGGCTGTACGAAAATCCCTATGTAACATCATCTGTAGATAAAAAATGTGGTTACAGCATTGAATTGTATCTAGATAACAAGTACAAAACACTAATGTTCTCCGATTTACAATTGAATGCTGACTATCCGTTGTATTACGATTCCTCACTGGATAAT tpg|BK006936.2|:718587-719809 7X164=1X186= 175=7X 
 tpg|BK006947.3| 107784 + tpg|BK006947.3| 108470 - INS CACCTTAAACTGGTGCTATGCATGCATGACGAGTCTGATATTCCGATTTTGTCGCAAGGGTTTGATGCTTTTGATGGATTGGTTAGGTCTGAATTTGTCCCTAAAGTAGTGGAAACGCTACTAAAATACCAAGATGACTTGATTAAAGAACACTCAAAGGATATACAAGTTTGATGTGTTCATGTAACGAAAAGGGGAGCGTTGCATAGAT tpg|BK006947.3|:107348-108906 28S84= 47=66S 
 tpg|BK006945.2| 345659 + tpg|BK006945.2| 345862 - INS GCTCTATTGACATGATGAATGAGACGATGAATTCCTTAAGATTTTGTTGTAGGCTTCGCTAAACTGGCTGATTCCATAATACATGTGCGAGAGTATATTCTTGTTATTATGTGCCTTCTCTCTAGTGTTTATTGCTACACTTTTATTGCTCTATAGTGCGTTGTATAAAGTAGCCACAATGGATTGTTGGCATTACTACAGCTTCATTATTTACTGAAATTTCTTAAAACGCGTTAGATGATATGTTGAAAAAAAAATACGCGTCGTGAATGAAACTTATTAGGTTTTACGACTAGTTAAAGCAAGAGAGAGAAGATCGAATTGACTAAATGTCTTCACTTTGAATTTATTCTAGTAGGATTCGCATGGCTTTTTCATAATAAAAATCTCGTTTATTTATGCTTTTGGTTGGTTTTCCTTTGATAAATGCGGCCCTTGCTTTGTTTGTGGTTGCAACGAGTTCGTCAAATGATAAATTGACGCTTAACACAGACGCATGGGAACCACGTAATTGAATTAATGTTTTCTTCTCGAAACAATTGCAATGTGACTTTCTTGTTAGGCAATGTGAGATGAAAGATGGCCTTTACCTTTGCAGATGTTTGGGTGTGGCTCTGAGCTGTCCTTTATAATTATAGAGATAATTTTGATGAAAGCTCAGAAGACCTTTAATGACGAAAAATAGGCATGGTTTGCCAGGCAAAAAACGACCAAATTTTACTGTAGTATGAGTCAAAGTC tpg|BK006945.2|:344165-347356 7X281= 370=7X 
 tpg|BK006936.2| 721845 + tpg|BK006936.2| 721956 - INS CGAGGCTTTCACGAAAGCTCAAAAGACATTGGATGAGGTTGCCCTGGGTAGAGGCAAAAAGCTTGTTGATGTCAGGAAAGTTTACTATTCAAGCTGAAATACTATGTACATACACACGCACCATTATCTCTCGTTTTACATAAGTAAATACAGCAATAATAATACCTGTAAATATCTCAACATAC tpg|BK006936.2|:721461-722340 7X124=37S 1S1=230S 
 tpg|BK006945.2| 875675 + tpg|BK006945.2| 875865 - INS CTATACATGATATATATAGTTATATATAGGTCGGAGCCAACAGAAAGAGCACCGATGGTAGCACCGCCGAAAGCAGCAGCAGTTGGAATGATCTTCTTCAATTCTCTGTAAATGGAGGTTTCTCTCTTACCGTTAATGACCATGCCTTGATCTTTGAATTGTTTGGCAATGTCACGTGGGGAAGTGCCGGAGATTTCGATCCATGTCTTGGAAAATACTGCGCATGAACCAAGAACAAATGTGATGTAGACGATGGTCTTGATAGGGTCCAGAAGAGCTTCGGATAAAGACATTAATGGTTGGATGTAGTAGACCAACCCGCTCAAGGCCATTTGAGGGCCCTGGGTGCCCGGCCTGATACCCCAAACACCGATCAAACGAATCAATGGATTGGTTGGGTATTTCTGGAAAAGGATTTGAGAGATCAAGAAAATGTTAGAAGTCAATGCACTCTGCAACATGATTGGGGTGTTGGAAGTATAAAAGAGTTTGATGGGGTAGATACCAATTTGACCTCTCACTTTGGTTGACC tpg|BK006945.2|:874597-876943 7X395= 10S286=1X219=7X 
 tpg|BK006947.3| 621699 + tpg|BK006947.3| 622268 - INS ACTTTGTTCCTCCTTCATATTTTTTTGGTCCTAACCTTCTTCCTGCAGAATCCTTCATACTTGTTCTCGAGCCCGCAGCCCTTTTGGTGGCATTACGCACTTGAAGGAACACACCAGACACATGTTTTTGGAATGAAAAACTAGAAGTATCTAGTAAAATAGGATTCCACATATTCTCACCTTAGGTTAAGCTTGAAATATTATGACCACCCAAACTGGCGAGTTTTATTTTTACAATGAGCCAACTTCATTCTTCAGTGAACTATCTTGAATGAGTCTCCAAAGAAAGAGCTTTAAAATTCAATAGCGGAACGTCAGATATCGAAACACCCAGTCATAACAGCCAAATTTGCATAATTGGTATAAAAACAGTGTGTATAAC tpg|BK006947.3|:620921-623046 7X250= 359=7X 
 tpg|BK006947.3| 181322 + tpg|BK006947.3| 181390 - INS TCTTGGACCTCTAGGTATATAACATTTCAGGTAGCTTAAATGGAACTTTCATAGTGGCAATTTTATAAGAAGCTGCAGTACTTTTTGGAATGCCAAAAGCCTCAGCTTGAGCCACTGTGGCACCTTTGACAATAGCACCAAGTACCCTGAACAAACTGACAACTTTGGAAGGTTTCAAGTTCAATTCGTGTGCTAAGGGTGTGATTTCAAC tpg|BK006947.3|:180886-181826 7X202= 185=7X 
 tpg|BK006947.3| 118527 + tpg|BK006947.3| 119114 - INS TGGTAGGGATGAAGAGAGCCACTAGAAGGTATCCCGACGTCGATTCCCGACGCTAGGTATAGGCATATGGCTCGATTTGAAGGACAGAATACCGTATTACAAGTCAGATTGGGTAGATGCGTTTAATTACAGAGTTATTCCCTCTATTGTTGACACCTACTTTAATAACCTGCTACCTGCAATAGCCTTTGCGCAAGATATGTTTGATAGGACTGATAATTCCTATGGTGTGAACGAAGTACTTCTATCCAGTGCAATGGCTGGAATTGTTTTTGGAGTTCTTGGTGGACAGCCCTTATG tpg|BK006947.3|:117913-119728 28S126= 150=7X 
 tpg|BK006945.2| 1007073 + tpg|BK006945.2| 1007674 - INS ATATATTGATGAGACAGCATTTGTTCAGGCTGAGCAAGGTAAAACCAATCTAATGTTCTCTGACGAAAAGCAACAGGCACGTTTTGAGCTCGGTGTTTCCATGGTTATTTATAAGTGGGATGCGTTGGATGTTGCCGTAGAAAACAGTTGGGGTGGTCCAGACTCAGCTGAGAAGAGAGACTGGATT tpg|BK006945.2|:1006685-1008062 7X6=87S 90S4=7X 
 tpg|BK006947.3| 208976 + tpg|BK006947.3| 209107 - INS GCCGAAGACTTGACCATCGCTGCGAAGACGCACATACTCAGAATTTCATTCTTGGATAGAAAAAGGGCCAAAGAATTTATTACGACTTTGTTGAAAAGCCTATACTCGTTTTTCAACATTTCTCCTGATGCGCCTAAAGAGATTATGGATAAAATAATAACAAGTAGGCCA tpg|BK006947.3|:208620-209463 7X4=246S 86=7X 
 tpg|BK006945.2| 125782 + tpg|BK006945.2| 126369 - INS TTTGGTGAAACGAGCTTTTTTGAGATAATGATGATTGTAAGAAACTTGTGCGTTGGTGAGAGCTTGTTCTCCTTTGTTTGTTACACCATCTTCAATTACCTGTTTGATTGGAACGATACCCTTTGGGATACCGCATTAAGAGATCGCCATTTCCTGTTTTCGCCAGTCCATGTTTCAGTGAAGTTGATGCAATGGTGGCTGTCACCCGACCCCAACAAGGTAAGTTTTAAATTTGGTTCCCATAAGATGTTCCCCGACAATGCTAAGTGGTTTTCAGACGCATCAAAGGCCCCAAAT tpg|BK006945.2|:125174-126977 7X148= 132S10=99S 
 tpg|BK006936.2| 746073 + tpg|BK006936.2| 745774 - INS CATGCTACATAGATTTCGTTCAAGCAGAGATATTAGATTGGACTAATCCTCACGATTTTATAGATAAATTTGGACATGAAAATGAATTTGACGTCATATTGATCGCCGACCCGATATATTCGCCTCAGCATCCGGAATGGGTAGTTAACATGATATCGAAGTTTTTGGCGGCATCAGGGACCTGTCACCTAGAAATACCTTTAAGGGCAAAATACGCCAAAGAACGAGAGGTTTTGAAATTATTACTAAAAGAGAGTGATTTAAAAGTAGTTGAAGAACGGCATTCAGAGGGTGTGGATGATTGGGGTGCCGTTAAGTATTTA tpg|BK006936.2|:745114-746733 7X8=169S 303=7X 
 tpg|BK006947.3| 468372 + tpg|BK006947.3| 469018 - INS GTTTGAAACAGATACTATCCTGAAGACCAAAAGCCCTTTCATAAAGGAAAATTTAAATGAACTTTTTGAAGCCGTTTTGATCTCATCTTTAACTTCTGGCGAGTTTAATAGATTATCACTTGATAACTTTGGTTGGGCAAGAAAGATTGTTAGATATTTACCGTTCAAATTAGATTCCCCAAATACTATAATGGCTATGATGTGGGAGTTTTTCTTACAAAAATATCTTCACAATGGTAATGCCAAGAATGATGCATTGTCTTTAGTTGCTACTGAATTCAACACTTACAAATCCACACCAAATCTTGATGAACAGTTTGTCGAATCCCATAGATTTCTTCTTGAAATTTCAAAAGTCATGCAGGAGCTAAATGCTGCGAAATTAATCGATGAAAACGTGTTTAAATTATGCACTAAAGCAGTTGAGTTTACTACAACAGCTCTATCTAGCTGAAGCGTGAGAATGAGTATGATGGAAATAGTGGAACTATTTAAAAAGCACCCAATAAAGAAAGAT tpg|BK006947.3|:467324-470066 7X279= 13S375=1X106=7X 
 tpg|BK006947.3| 474099 + tpg|BK006947.3| 473547 - INS GGGCTATATCCTGAATCTATCGAATGTTCTGATAATGGTGATGGCATAGACCCTTCAAATTATGAGTTCTTAGCTTTAAAACATTACACATCAAAAATTGCGAAATTTCAAGATGTTGCTAAAGTACAGACGTTAGGGTTTAGAGGGGAGGCCCTATCTTCTTTATGTGGCATAGCTAAACTAAGTGTGATAACAACAACTTCACCACCAAAAGCGGATAAGTTGGAGTATGATAT tpg|BK006947.3|:473061-474585 7X4=5S 222=7X 
 tpg|BK006945.2| 146863 + tpg|BK006945.2| 147435 - INS AAAGAAATATTTACCTCAGAATGGCAACAAATCTTCAATCTTTAACAGGGAAGAGGGAGCATCGGGAGAGAAATCAGCCGGTTCCTGCAAGCAACATCAACACGTTGGCGATAACAATGCTAAAACCGCGTAAAAAAGCTAAAGCCTTGCCTAAAACTTGATACATATTGATATTTATTATTTAGTACACGTATGTAGCATCGATCTTAGAAAATGCATGTTTGTATTTATTGTTAGTACCTTGATCGCCACCTTTCTAGGTAATGATAGGTCCTCAACTTTTACTACGCGGTGCACGCCTGTAAGG tpg|BK006945.2|:146235-148063 137S233= 288=7X 
 tpg|BK006947.3| 77041 + tpg|BK006947.3| 77215 - INS GTGCAGGAACTCAGGTTTTCCGTCTGATGCAAGAAAGGGTAAAAACTTTCATGAGTTAGACGACGTTCTTCCCAATATACAGGTAGTGGACGCTTCCGAGAAAGATGGCAAACTCAATGTGCAGGAGATTATTGAGGACTTACAAAGAACAAGTTTGAGAGAAAGCATTCATAGTATGGAACAGTTACCATCTTCGCACAAACGTAAACCCGTAATACCGTGGGAC tpg|BK006947.3|:76575-77681 7X4=123S 113=7X 
 tpg|BK006936.2| 579586 + tpg|BK006936.2| 580102 - INS CCGTATAGGTGTTTGTCTTAAAGCTTCTTTTTCCTTTTGTTCCTTTTGTTCCTTTTGTTTCTTCAATAAATCATCCTCTTTTTGCTTTTGTTTCTTCGATAAGCGAGCTTCTTCCTTCCTTTTGAGTTCTCTGTTCCGTTTCTCTTGTTCATCCAATAACGCTTTTGCTACAGATTCGGATTTTTCCTTCTTCCCTTTTTCCAGCATAGTGGTCGATTTGTATTCTTGCTTGTGAGATTCATCTGTTTGACTAATGGTGGTTGCTGAGGCTAATTTAATATCGACTCCCTTGGAGGTGGTACCTCCATCCATATCCCAGATATTGTCATGTGTCAATGGCTTGAAAATATCGTTTTCAGTAGCTTTAATAGTGCCAGTAGCGGCAACACCGCTTGCGTAAGGAGCTAGATTCAAGTTGATAGAATCAGAGCTGGTTGTTTGAACGTGAAGTTTGTCAAAAGTAGTGAATGGATCCGTATCATACTTCTCGAGTTTAGTCATTAACTCACCAAGTGTGATGAAAATATCGTTTATTCCTAGCGTTTCTGGAG tpg|BK006936.2|:578470-581218 7X134= 2S532=7X 
 tpg|BK006947.3| 239688 + tpg|BK006947.3| 239527 - INS CTGAGATTGTATGTTGCCCGAAGAATGATTCGAATAGCTTCTGAAGATATCGGATTACGGGATAGTTCATTATTGCCCTTGGCTGTCGCGGCACATGACGCAGTAATGAAAGTTGGTTTGCCAGAGGCAGACCTTGCACTGGCGCAATGTTGTGTTGCTTTGGCTAGGGCACCAAAGTCAGTAGAACTATATAGAGCTTGGAAGAAATTAAGGGCAATGATGAGCGAGAACATGTACAGTTTAGCAAGCACTGAGATACCGATGCATATCAGAAA tpg|BK006947.3|:238963-240252 7X233= 113=1X24=7X 
 tpg|BK006945.2| 164133 + tpg|BK006945.2| 164205 - INS AATGATTATGCAGTTTTGCAATCGATAGTACTTCCGGAGAGTAACAGGTTTTTCGTATATGTTAACTTAGCATCAACAGAAGAGACTAAGTTAGCCACAAGGTTTAACCAAAACGAGATCGAGTTTATGAAATGGGCCATAGAACAATTCATGATCAGTGGAGAGACTATCGTTGAAGGG tpg|BK006945.2|:163759-164579 7X5=85S 85S5=7X 
 tpg|BK006945.2| 798656 + tpg|BK006945.2| 799253 - INS CTTTATCTCCTTTCTTTCCTGCAAGGAAATTATGGTATCTAAATTTCTTGTTAATAAACCACTTCAAACCTTTGAGAATGAATAGCATATTTTCCGATTTAACGTTCTTCGTTAAAACATCGCGCAAATAATCATCGGAGTAGATTATACGCTTATTTCCACTTTCATCCATCTTGAGTTTCTTCTCACTTTTTTTAGCTACAGTTAAAAAT tpg|BK006945.2|:798218-799691 7X6=100S 93S9=1X3=7X 
 tpg|BK006936.2| 108615 + tpg|BK006936.2| 108404 - INS CTATTAAGGGATCGCAAAGAGGTATGTGCGCCAGTTTAAACGAGGTAAAAAAGAATGACACCTATGGGGTCTCACAAAAGGGCTACAATGACAATTTCAGTGAAAGTGAGGGCGTCCTTCATGGTAGTAAGTCGATGCCCACTAGCATGAAAA tpg|BK006936.2|:108084-108935 7X6=70S 71S6=7X 
 tpg|BK006947.3| 754672 + tpg|BK006947.3| 755166 - INS GCATTTAAAGAATGAGAATCTCTAAGGGATCATAGTCTAGAATGGTATTCTGCAAAACAAATTTTAAATGGTGAAAACTTTTCCTCACTATGTCCAATTGATGCTTCTTAGGATGACGTTAGAATTTTATTTTAGTGCAGGCATTACCTTGCTAAGTTCATTCATTAAAGTACTAATATACCTCTTACTGGCATGCATTTACC tpg|BK006947.3|:754252-755586 9S169=12S 14S6=7X 
 tpg|BK006945.2| 1011432 + tpg|BK006945.2| 1012156 - INS AAGCAGCATAGGTGATGTACTCCGCCCACAACTACCACCCCTTGCCCGTCGTTTTTCACAAGGCTAAGGGCGCACATGTGTGGGACCCGGAGGGTAAGCTGTACCTCGACTTCCTGAGCGCTTATTCTGCCGTCAACCAGGGCCATTGCCATCCTCACATCATCAAGGCTTTGACGGAGCAAGCACAAACACTAACATTGTCCTCCAGAGCGTTCCACAACGATGTTTACGCGCAATTCGCCAAGTTCGTGACCGAATTC tpg|BK006945.2|:1010898-1012690 24S113= 26=111S 
 tpg|BK006945.2| 1014566 + tpg|BK006945.2| 1014922 - INS CGTTCATCTTATTCACTTCCGACTTCGAACCTCATGCCGTTCAAGATGCTTGTGTCGCCATCAAAGACCTGAGAAAGTCCCCAGATAATAAAGTCCCTAAATTAGACGAACTCCCCACCGTGAGAAAATACTTGAAACAGCTAATTCATGCAAGCTCCGTGGAGCAAGCAACTGCATGATTCCCGTGGGCTTCCTACCCTCTCTCCTGTAAATATATATATATATATATATCCACACACACTCGCACATACATACACACATACATACACCTTTATATAGCTATACGC tpg|BK006945.2|:1013978-1015510 7X46=1X192=21S 3S1=449S 
 tpg|BK006947.3| 606054 + tpg|BK006947.3| 605335 - INS GCCCAAAAAATATATATACAAACAAAAAACAAGGTCCATAATGACAAAGAATTTCATCGTCACTTTGAAAAAGAACACTCCAGATGTGGAAGCTAAGAAGTTCTTGGATTCAGTTCATCACGCAGGTGGCTCTATTGTACACGAATTCGACATCATTAAAGGGTACACCATCAAGGTACCAGATGTTCTCCACTTGAACAAGTTGAAGG tpg|BK006947.3|:604903-606486 7X6=154S 183=7X 
 tpg|BK006936.2| 783364 + tpg|BK006936.2| 784007 - INS TGAATTCGATGATATATTGTAACGGCTTGGTTTGCGGCCTGTCTCATGGAAACTGGCAAAACACCACGATAAAGACCAGAAAATCCTTTATCACGGACTAATGATGAATAGTTTCGTACTACACCGCGCCCATTATTATGGTATTTTGGTGTAGCAGATTGTTTATCATCGATCAAAGCAGTTTTGATTGCTTCAAAAGGAGTCACTGCGGCAACACTTTCTAATAGTCCCGCACCTAACCCAGCTATCACCCCTCTTGTACCACTTAGTTCTCCAGTTTCACTATCTCTTAGCATGTCTTTAATGG tpg|BK006936.2|:782736-784635 61S207= 288=7X 
 tpg|BK006947.3| 79621 + tpg|BK006947.3| 78890 - INS CTTATCCACTATTATTGTGGCCTACGCTTTTCTGGACGATTTGGTCTGTAAAGTATAAAATTTTATCACGCGCATAGCCTAATTTCTTCAGCGCTACATCTTTATAAGTTCCCCTATCATTGAAATGCATTCGATCAATGCTTCTGCCCACTGATATCTGATCTTCTGGGTCGTAGCGTGATATGGTCTGTAAATCACATACTTCCGAATTACTTGACGTATCGTGCCGATCCGTTGATGCGTCCTGAGATTCCCTCCTGGTTAAAGCGTTTTGAACCCTTAAGGCGTACTTGGCAAACCGATAGTCTTGTTGCTCTTCCTCGAAGATAGGTCTTCCCAAAATGCTTTGCGCTTCCTCTTTTC tpg|BK006947.3|:78150-80361 7X8=172S 341=7X 
 tpg|BK006936.2| 548039 + tpg|BK006936.2| 547851 - INS ACTACGAAATTGGAAGAATTCTTATAATAACTATTGGATCAACATTTCTGGGTAGCTCAGGCACCGAAGTTAGCCCACCCCAAACAGTAAATTTAAAGGATATGTCATGGTGGAAGGGCATTACCGATGTGGTGCTTTGTGCGAGACTGGCCGATGACTAATAGTGTTAGAACTCCACCTTCTGTGTAATTTCTTTCTGAAATTAGTGAAAAAAACGCGCCTTTCAAATTTTCATACTAGTGATTGGTTTATTGCAGATTATTTATTTCTAATTGTACATATTCTTGTTATTTTATATTATATGAAAGGGGTAAATCCAAATGCCACTCTACATACAGATTCTGTAACTGGCATAACGACCAGAGG tpg|BK006936.2|:547105-548785 7X137= 344=7X 
 tpg|BK006945.2| 352957 + tpg|BK006945.2| 352857 - INS GTTCTGAAGTTGCTGAGTATTTCGAAATAACAGACAAGGTCTGTGCGGCATAGTCTAACAAAGAAGGCAGCCACTTTTCAAACAATCTGACATTATCTACATTCGCTTTTAATGAAGAATGAACAATATCGCCCTTTAAGCAAGTAAAGTGTTCTAGGTCTAACATCATACCATTAATCTTACAGTAATCATTCGTGAACT tpg|BK006945.2|:352441-353373 7X5=95S 88S13=7X 
 tpg|BK006947.3| 576212 + tpg|BK006947.3| 576755 - INS GTAACACGCTTAGCGTGAATAGCAGCCAGATTAGTGTCTTCAAACAAAGAGACTAAGTATGCTTCGACGGATTCTTGCAAAGCACCGATAGCAGAAGATTGAAATCTCAAGTCGGTCTTGAAATCTTGAGCGATTTCTCTGACCAATCTTTGGAAAGGTAA tpg|BK006947.3|:575876-577091 7X4=76S 75S6=7X 
 tpg|BK006936.2| 656465 + tpg|BK006936.2| 656626 - INS TATATACCATTCTTCCTCCATTATAGGGGGAATATAGTTCCTGCAGAATGTGTACACCCTACGAAGAAGGAAAAGGGCATCTTCAAAAGTGTCCGCATGACTATACACAAATTTCTCAATTGTTGACACAGCAGCTCCCAGATATTTCGAAGGAAACAGAGTAGAAATCCTTTTCAGACTCGCCCCTATGAATTCAAATAAAATGTAGGATTTCAACTTCAAGAAAAATTCATTTGAACTCTTGCTTTCACCGTAGGATGGAAAATCTTTTCGATTAGAGGAATTTTCGATTACTCCTTCAGGAGGTAACGTATTGGCCTTTTTATCAACAAAGTCTTCCTTATTCTGT tpg|BK006936.2|:655753-657338 7X171= 3S325=7X 
 tpg|BK006936.2| 727931 + tpg|BK006936.2| 728319 - INS AGTTATACCTTTGCATGTCACGTGAACCAACAGAACATGGTAATACATAATGAAGAGAAGTTGCCTAAGTACCTTAGCTACAGTACCAAGTTCTAATCTCATCATTATCACACATTTACAAGACTATTTTTGCAGCAGATGGAGAGATCACTTCAAAAATGCGTTTATGAAACCTATTTATGACGAATTTTTTATTTATTTATTTAGGTAGTTTCTAACCTTCTCCTCGATAATGTTTGAGATCATAGTATTCAAAGTACTATCTTTCTTTGATATTTGGTTTTCCAACGTTAATAGAATTTGCTTCTCAATAATCTTCCCAGTCAAATCTACTTCAATATTAACCTCGTCGCCAATTTT tpg|BK006936.2|:727197-729053 7X4=209S 180=7X 
 tpg|BK006945.2| 98532 + tpg|BK006945.2| 98989 - INS CCTTTCGTCTTGAATCTGTGCGAGCCTTGCCTGCTGTAACTCGCTGTCCTTGGGTCTTGTAGTCATGTGTTTTTCAAGCAGAGCCTTGGCATGCTTGAATCTTTTTAGTTTGTCCTTAGCCGGCACCTGATCAACCCACCTTAAAGCATCACACACCAAAAATTCTGCTTGTATCACCTTCTCAGTTACTTGTTCTGCGGGTTTCAAGGTCTTGTAATAGCCAAGCGCCTTCAAGTAATGATGAATGGCTCTACTGAACATCTCCGCCTCCCTTTCGATGTCACCCATCAGGATATACACATCACCGATGCGCAATCTGCTGTTCTCGGTTAGAGATTGGCCATCTGCTGTAGGGCGGCCCAACAGCATCAAGGCCTGCGCCAGTAGGTCCAAAGC tpg|BK006945.2|:97726-99795 7X157= 198=7X 
 tpg|BK006945.2| 855801 + tpg|BK006945.2| 855689 - INS CCTCAGTTGTGTGGTTCAAAGTATGTGGATCTCCGTCTCCATATTTCAAAGGGAAGAGAACAATTTGTGAACAAATAAATTATAAGATACCACATTAACAACAAGTATGTGGACGAGGTGTGGTAAGATCTCCGCTGAGGTTGATTGAAAAGTATTGGGTAAATTTGTACTTTTTGTCTGCTGCTGGTCGTTTGTCTTTCGTTTTAAAATTGCGCTAGACAAGTAAACAGGGATTGCTTAAGAATCAAAGTAGCTTAACTCTAAAGTATTATTTTCCTCAGTTGTGGGCCCATGTGTTGGAG tpg|BK006945.2|:855071-856419 7X266= 29S236=7X 
 tpg|BK006936.2| 210392 + tpg|BK006936.2| 210785 - INS GTTTGAGAGAAATAGTAAAAGGATTGAAAATAATGTAAAATCATCCACCAAGACCATTAACAGTAAAAATACATTGCTAAATGTGCCAGAAGGCGTTGAAAAGAAAATTAGTATCTCATCGTTCCCATTGCCAAGGTTGGGCATACATTCTTTGATTATGGGTACAAAAGAAAGGAGTGCATGGAAAATCTCAAATTCAGAGCTGGAGAATGATGATGCAGATAATGCGGGTGGTAAGGGTTCAGATGGTACGAGCAACAGTATTGACGACATTGCAGTTCTCTCAGAGGAAGAAAATGACTTTCATAGGATGACTTTGAACGCCAAGCTAACCCAGGAGAAGAT tpg|BK006936.2|:209688-211489 18S161= 121=59S 
 tpg|BK006947.3| 417128 + tpg|BK006947.3| 417502 - INS CTCTCACTACTATCGCTTTTTGGCCACGAATGCGACAAAAATTTTCTCGTTATGCTAACCTCTCTCACTATCTCGATCTCGTATAGCTTTCTTTTTTGCAGCTATTGTTCTTTTTCTGGGCCGTTAAATTTTTCATCCGGAAACTCCAGGCTATTACCCGCTCCGTGATTTTGGTCGTTGAATCTTCGTAAAAGCAATCATGTAAATATCATTGAATACGGACAAACGGAACTATATTGCTGGAATTAATGATATAAATGGTTTCCCAAGTTTGCTATATCTCCTATTC tpg|BK006947.3|:416536-418094 7X393= 271=7X 
 tpg|BK006945.2| 330620 + tpg|BK006945.2| 331112 - INS CAGGGACGTGTAGTGGCTTTCGAACTTTTATTCTCTGACCAGTATTCTAGCATGGACCCCCAATTAGTTGTAATCACATCATAATCAATTGTAATCGATTGAAGATATGCATCGATATCGTGAGAGTACTCGAGATGAATAAGCTCCACTGAATCAGGAATGTCTGGGTCGCTTTCTTTTATAGTACAGTTCTGTAGTTTTATTGGGATATTCAGAGTTTGAGAGACTTGGGAGGAAGAGCCTTCTTTTACTCTGTGAATGGTTTTCTTTACGAGTACACCAACATTGGGTAAGGCAAACAAGCTCTTCATTTCCTCCCCTCCACTATTATCATCATCCAGTATAACTTCACTAAACGTAAACAGATGCAAGTTATTCGCTAAGTAGTTTTTGAAGATCATATTTTTCATTTCAATTAATTTTATGATACTGTAAATGATGTCGAATTGGCGTGCAATTTCAAGC tpg|BK006945.2|:329676-332056 7X228= 451=7X 
 tpg|BK006947.3| 171120 + tpg|BK006947.3| 171273 - INS TTCCAGCCAAAATGTGTGACTTCACAATAAACTCAGCAGTCCTATTTCTCTCGTCCTGCAAAACACCTATGGGCGTAGCAGAAACAGACCAAGTGTATATCTGATCACCGCTCAACAATTTCAATTCGTTCTCTGCGTGTACGTGTAACGGCTTAGATTCATCAGAAAGATCGAAGTTAGGGAATTTCCAAGTACCGCTT tpg|BK006947.3|:170706-171687 7X119=31S 2S1=78S 
 tpg|BK006945.2| 872998 + tpg|BK006945.2| 872953 - INS ATAAATACCATGCAAGATTAATCCCGTGATGTTTATGCAAGATAGCGAATTCATGTAGATCGCGCCATGCTGTCTTTGCTTTTGTTGGGACCATATTGATACTATATCTATGATTAGGATCTTTTCGTCCCCCGTAGTACAATTCACCAACTTTTGCAGCGCTACCGAAGGTTTAAAATCACTTTCAATGATGTGCAAGAACCCTAGTTTACTCTCCTGCTCTTCACTAATTAGGTTTCTTAATTCATTTGGTAGGTTTATATAGTTCTTGGTTGATGTGATGAAGTTTGACAAAGGATAAATTCTAATGTTCTTTAAAACTTCCATCCCATTCCATTCGCTACTTCCTTTCTCTTTTCCTAAGAATTTTCATTATTAGAAGGAGTAATGCTTACGGTACACATACATACACATATATATATATAAATATATATATAT tpg|BK006945.2|:872063-873888 7X116=1X191= 2S423=7X 
 tpg|BK006945.2| 952185 + tpg|BK006945.2| 952434 - INS GACAATTACGATGTCATTATTTCTGGCTCTTCTCCATTTTATGGCCTAATGTGGTCTGGATTTGTATTTGCCGTCCTTGTATTTCTCTGCATTGCATACTGCTGGTGGAGCAGCAGAAAGGGAGCTGCCATCGTGGAAGCTGAGAAAGCTGTTCAAGAAAGTGACTCTACTACCTCAAGAATCATTGAAGAACACGAAAGCCCCATTGATGCTGAAAAAAACTTTGCAAGGTAAAATAA tpg|BK006945.2|:951693-952926 7X5=114S 114S6=7X 
 tpg|BK006945.2| 949781 + tpg|BK006945.2| 949704 - INS GCCCTCGAACAATACAATATTGTTCTTGATTAATGCATTCAAATATGTAACTTCGGCCCTCATATAAGCGTCTGACGCGTCGTGAAAATTTACCCTCGCAAGAAAATACAAGAGATTACGTAAAATTAGAAACCAAAAGATATGAGTGGAACAGACACATATCACCCATATTTCCTTTTCACGTAAGAAAACTTAAGTACTAGTGCGGTGCCTGCGTTAGTGCTTGTCTTTAGGTCAAACAGGTCATCTTGACC tpg|BK006945.2|:949182-950303 7X412= 40=1X41=1X156=7X 
 tpg|BK006947.3| 481418 + tpg|BK006947.3| 481301 - INS GATTATAATACAGTGATAAAAACAATCATACAGAAGAATCCAAGCGAAAGTTTCAAGAGATATGCCAGGCATACGAAATACTTAAAGACAATCGTTTAAGAGCTTTGTATGACCAGTACGGTACCACAGATGAAGTCCTGATTCAAGAGCAGCAGGCGCAGGCGCAACGCCAACAAGCCGGGCCGTTCAGTTCATCCTCAAATTTCGATACGGAAGCAATGTCATTCCCGGATCTATCTCCAGGTGATCTTTTCGCGCAGTTTTTTAATAGTTCTGCTACCCCC tpg|BK006947.3|:480719-482000 7X6=147S 267=7X 
 tpg|BK006947.3| 435997 + tpg|BK006947.3| 435943 - INS ACCTTTATCTTATTTTTACAGCCAAAAGGTTGTTTTTTGACCTGATGGGGACCCCAGCAATGGGTGTCGTCTATGGCTTAAATGCAGACCGTTGGACGCTGTTTATCGGGACGGCAATATTTGCTTTCGAAGGAATCGGGTTAATTATTCCTGTTCAAGACTCAATGAGAAATCCTGAAAAATTTCCTTTAGTACTTGCTTTGGTGATTCTAACGGCAACCATACTTTTCATTTCCATAGCTACATTGGGATATTTGGCATACGGCTCAAATGTTCAAACGGTTATACTGT tpg|BK006947.3|:435347-436593 16S136= 93=60S 
 tpg|BK006947.3| 712064 + tpg|BK006947.3| 712774 - INS GACCCTTTAAGGATGAGTAGTGTCGTTAGTATTCCATTGAGAGAAATTTTATGATTGATTATCATTTACTATAAAATCCCTGCGTTTGATTCGGTCTCTAGGGAAGCGTTGTAATTTCATGTATATTCAAAATAAGGACGAGGTTATATACCATACTATATTATCTCCTTGCATTCTGTATCAAACACTTTATTCAGTACATATACGATACCTATATATTCATTAAATGTTCTTTTCGCTTTATTTCAGCAAGGTATAGTGCTATTTAAAATCCATAATCGTTATTGCGTCTCTTTAGTCTGTCCTTCATTGCCATTACTCCACTACTTGCGTCTGGTGGCGGCGTTGGCGTGCTGGAGGTGTTGAAACTG tpg|BK006947.3|:711308-713530 7X299= 348=7X 
 tpg|BK006936.2| 137086 + tpg|BK006936.2| 136909 - INS GACTACGACAGAGGAAGAACAGGACACTGAAACGCTCGATGCTGTGAGTTTGCATAGTTCAGCGCCAATCTTCCGTGTGCTCTCTCGGCGGGTAAATGGACAAGAAGATGACAGCGAAAACGAGAGTAGTAGCGATGTCGACGATGGTTCCGTACCATTAACGAGATTTCATTCTTGTCCTATCACAGCATAAATTAAAATGAAGGAAATAACACAACTTCGTTTTGCATTATCATATTCACATC tpg|BK006936.2|:136405-137590 7X263= 123=7X 
 tpg|BK006947.3| 378135 + tpg|BK006947.3| 378232 - INS AATCAACTCCACTCCGTGTCGAGCGGTTCTGAAGCCGTTCAGGCGATGAGGGAAAAACAAAAAGAGCTAATCAACTCCTTGAACTTAGATAAATACGCCATAAATGATAACAGTGAGGAATGGGCTGAATCTCAAAAATCTTTAGAAATAGCTGCCAAGGCCAAAGGCGTCGTCAGTTTAAAAACTGGTAAAAAGAGAACGACTGAAAAGGCTGAAGATATCTATAGACAAGAGATGAAAGCTATGAAAAAACCAAGAAAGTCTAAAAAGGCTGCAAATTAAGCGTTCTACTCTTTGTCAAACCCTTTTATAGC tpg|BK006947.3|:377493-378874 7X8=223S 4S291=7X 
 tpg|BK006936.2| 541088 + tpg|BK006936.2| 541622 - INS TCTTCATTGTCAAGGGCATAGAATTTTGCGTATTTACTTGTCAGATTGAACTTTTCCATCGTACTCCGTAGAAAAAAAGTGTAAAAAAAAAGAGATGTTTGCCACTTCAGATTGTGTACTGAAAGACAGCGTTCTTCAGATCCAAGCATACGGGTATGTGTATCCCTCAATAATCCAATTATATAACCAGTCTCCATGGCATGTTCGTCATTAACCATAATCTCTGACAAATAC tpg|BK006936.2|:540606-542104 21S103= 31=93S 
 tpg|BK006945.2| 143515 + tpg|BK006945.2| 143754 - INS GTATGTGAATTAAATATTCGCAACAAATTCATTGCATTGTCCCTTGCAGAATATACCTACGCTAAGAACAAAATCAGAAGACATTTTAATCACTGGAAGACTGTATGTGAATTGAATGAAGAGGCAAACAGGTTTGCAAATCAAGCAAAGCGGAGGGTACAGGAAGCCGTCTTCTATATTTGGAGTGATAAAACATTAAAATACTCACAGATGGCCAACGATGAAGCTGAAAGTTTTAGGAATACTTGGCTACTATTTCGCTCGTTCCAACAATGGATAACTTTAACACAAACTCTTAAGGAGCAGTCAAGGTTAGCAGATCAGGCCTTTTTGAATAAGATGTTTAGGAAAATTTTAAAGGCACAAGAGCATTGGAAACACTTAGAAACTGTTAACACTGACAACATTAAGAAGATATTTTTACGAACAACATTTCATATATGGAAGCTAAGACATAAAGAAATAAAC tpg|BK006945.2|:142565-144704 7X325= 3S134=1X316=7X 
 tpg|BK006936.2| 144371 + tpg|BK006936.2| 145132 - INS AACGTGCGAGTATATTTTACCAGTAGTAATGTTATGATCTTTAGTCAAAGTAACTCCAAGGTATCTCTCGTAGTTACCCAAGTCCAAATCTGTTTCACCACCGTCGTCAAGCACGAAACATTCACCATGTTCCAAAGGAGACATAGTACCTGCATCAA tpg|BK006936.2|:144041-145462 7X25=54S 1=200S 
 tpg|BK006945.2| 65633 + tpg|BK006945.2| 65219 - INS CCTCTGGTGGTGGGATACCGGTCAAAGTAAAGTGGGAGGGAGAGTTCGAGAGTTCTTGTCGTATTGTAGTAGATAGAAGATATACTTATCCTTATCCGTACAGTTCTTGCTCTTTCTGAAGTAGCACTTTCGGAAGAAGAAAGATAAGCAGGCGAATTCAAAGGTGGCAAAACCCGGAGCCTCTCTATATATACCCCCAAAAGGAGGAACCGCCCTCAAATGACACTGAATTCTAAAAACAACTGATAAGTGGCATCGCCCCTGAAAAAAGAAACGAAGTGGGGTAACCACCGTGTGTGGCCGGATGTACGGCTGTGTGATGCTCCACTGGGCGGCTATTTTTTTTTTTGGTACCGAAATTGGTTTATCCAGGATTATTCTAGAACGTTCTAGAAACAATACTGACCACAAAGACTTTTCGGAATAGAATATTGTCAAACAAGAACTTTTTCACTTTCTTTTCATAAAACGTCACTTTCATCACTTTTGCAGGATTTCCCACAGTTCGTTTAAAGGGACATTTCCTATCATGGGTTGCCCTGCGCGAATAAGATGATTGGTCAAGGAAGACTCTAAAATCATCTGAACGGGTTATTTGAAGACTTGGGTCTAAATGAGAGCTTGCTTATTCCACCCGCCACGCCGGGCGTATC tpg|BK006945.2|:63899-66953 7X4=172S 3S630=7X 
 tpg|BK006947.3| 710015 + tpg|BK006947.3| 710186 - INS AGAACCTAGGAGAAAATAAGATACCATTCGTCATCGTCACACTATACCATTCGTTCCAATCTGAAGACTATTTGTATCTCTGTATGGAATACTGTATGGGCGGGGAGTTTTTCAGAGCTTTACAAACAAGGAAAACCAAATGTATATGTGAAGACGATGCCAGGTTTTATGCCAGTGAAGTGACAGCAGCACTAGAATATTTACATCTGTTGGGTTTTATCTATAGAGATTTAAAACCAGAGAATATTTTGCTGCATCAATCAGGCCATATCATGCTTTCTGACTTCGACTTGTCTATTCAGGCTAAAGATTCCAAGGTTCCTGTTGTCAAGGGTTCCGCTCAATCAACCCTTGTTGATACCAAAATATGCTCAGATGGGTTTAGAAC tpg|BK006947.3|:709225-710976 7X190= 6S358=7X 
 tpg|BK006947.3| 463070 + tpg|BK006947.3| 462355 - INS GAAATAGCCTTTGACTTTTTGTTCTTTAACGAATATCATTAAAAAAAAAGGACATCTATAAAGAATGTCTCCAAACTCGTCGAAAACTCGAACGGACCAGATAAGCTCCATGCCTGGTATTAATGAAGCCACGAAGGTGGAAAGTAAGAATGTTGTGAAGGATGCTGT tpg|BK006947.3|:462005-463420 7X12=147S 147=7X 
 tpg|BK006936.2| 181206 + tpg|BK006936.2| 181903 - INS CAAGGTCTTAGCGTGGAAATTTGCTGCAAACTGCCGCTGGAGCTAGCGTTTCCACCGTTCTCCTGAGTATCCTCTGGGCTTGTGCTAACATGTTCGGACTCGTTGGTATTCATATTCTCGAGAGGTTTGTGCCACTTGTGTTACTATCTAGCTTAGTCCTGCTCTTGAGTTTGATTGGCGGAAAGCTACTATTCGCAGCTCTTTTTTTACTTAGTCTGAAAGAGCGGACCAAAAAACGCACGTAGCGCGATATTGTCGTGGCATCGAACGTAATAT tpg|BK006936.2|:180640-182469 174S114= 138=7X 
 tpg|BK006947.3| 156003 + tpg|BK006947.3| 156040 - INS GTGGCGAAGAAAGAAGAAAGAAGTTAACCCTAGATATTTACAGCCTTCTTTATTTGCTATTGAAAGACTTTTGGCTATTTTCCAAGCTATATTCCCTATTCAAGGTAAGGCGGAGAGTGGTTCCCTATCTGCACTTCGTGAGGAATCCTTAATGAAAGCGAATATCGAGGTTTTTCAAAATTTATCCGAATTGCAT tpg|BK006947.3|:155597-156446 7X5=148S 98=7X 
 tpg|BK006936.2| 48676 + tpg|BK006936.2| 49162 - INS TTGAAGAGCTTCTATCTGACTCTTGCTGCAGAATCATTTAAGAGATTAAACAGGATCATGTTTGAGAACAATATTCCCGGAGATAAAAGAAGTCAACGGTTTTACATGAAGCCGGGGAAAGTGGCTGAATTGAAGAGATCTCAAAGGCATAGGAAGGAATTCATGATGGGCTTCAAGAGGTTGATTGAAATTGTTAAAGATGCCAAGAGGAAAGGATACTAATCGTACCATCAACTCTTGAATATTGTGAAATTTTCGCCATTGATTTCCGTCTTTGTAAATAGGTAATGCGTAACTATTTAGTTAAATTTTTGTATATTTTTTATTCTATGACTTCACTTATCCATTATTTCCATCGTCAAAAAAAGGAAATAAATACTGTTGCTCGAACGAACAGCAAGATAAAGTGGAAACGAAAAGTAAGCAGCTTCCTCAATATGCCGTCAAACGTACGTTCGGGAGTCTTAACTT tpg|BK006936.2|:47720-50118 7X153= 11S446=7X 
 tpg|BK006936.2| 344637 + tpg|BK006936.2| 345297 - INS AGTATTGCATTCAGATCATACTCGCCACTTTCTCTTAACCATTCTAATATAGCGTAAACGATGGCTTGACAGGTTAAAGTTGAATTGGGCGCATCATTTAGAGCCTCTGCACGTTTCAACCATGCTGACAAGGTCGCTTTGTACCCATTTTTAGAGAGTTCCAATAAACCCTCCTTGAGCAAACTAACTAGTTTATCTACAGG tpg|BK006936.2|:344217-345717 7X11=90S 98S4=7X 
 tpg|BK006947.3| 471290 + tpg|BK006947.3| 471506 - INS TTCTTGAGTTTTCTTGAATGGGCGTTTCCAAAGAGAAAAGCCAACATTGCGCTACGAGGCCAGGCTAGCCACAAAAAGAATACTGATAATGATCGGTCAAAGAAAACCACCGACTCAGATTTATACGTTACATATGATCAATGGAGAGACTTTTTGCTGCTGGTACCGAGAAAGCAGGGTTCGAGACTTCATACTGCTTATTCCTATTT tpg|BK006947.3|:470858-471938 7X4=1X3=1X3=1X150=19S 5S1=214S 
 tpg|BK006947.3| 16489 + tpg|BK006947.3| 16852 - INS CACTCGGTGGATAAGGCAACTGCGTATAATTTGTAGCTTCTTTTCAAAATATAGTAAATGGATATTAACATAAAATAATCACTTTAACTAATTGTCAAAAGCTATCCTGGCAGACATCGATGTGAGGGGTGAAAGC tpg|BK006947.3|:16203-17138 7X5=63S 62S6=7X 
 tpg|BK006947.3| 137519 + tpg|BK006947.3| 137670 - INS ACACAACACAGAATGAGAAAATGATAAAACCGAGCAACGCGATGACCTTTATGGAGGCAATACAAAACTCAAATTCTCCGTAATACTTTACGGGAAACATGTTCATTGAAGTTAACAGGCACCAAAAGATCACGATCCAAGCCGCTAGAGGCACTGCTTCTGTCCAGTACTGAATAACTTTCCCCAAAACGGATAGTTCCAGTGCGAAGGTGAAACACCACGACAGCCAGTACATATATCCGTTAGTCGCTCCCAGCGCTGGCGACAGAA tpg|BK006947.3|:136965-138224 7X3=176S 135=7X 
 tpg|BK006947.3| 769401 + tpg|BK006947.3| 769351 - INS TGTGGTGAATAACAAGTAAATTTAAGAGAAAATGAAGAAAAAAATTGCAGGTATACTATGGGTGCAGGTGAGGCGGTTTTTTAACCGATTTAGCACACGATACTGTGAATTTTGGGTTATATGATGATGTGAATATTGCAGAAATGTAATGTTATATTATTCAAAGAAATAGGGTAACTTCTATTTATGCAAACATTGGTAATCAAGGCTATAAACACATAATCCCAAAT tpg|BK006947.3|:768877-769875 7X6=1X190= 115=7X 
 tpg|BK006945.2| 518135 + tpg|BK006945.2| 518708 - INS TTATACAACGACATTGTAAAATTTAGCATATAAATTTTGGCTTTTTCTTGATCATGTATTAGCGTGTTCATAACGTGTAAGCTTTTGTCACTGTCTTCTGCTTCACTCTCGCCGCCAATCTCCTTCTTAAACGCTTCAATAGTATCAAGAAGTTCTGTCGCTAGTGCGGTCATCTCTTGCGACCGATCTTCTTCACTCAGTATCAATTCCACCGCATATAA tpg|BK006945.2|:517679-519164 7X5=105S 106S5=7X 
 tpg|BK006945.2| 832033 + tpg|BK006945.2| 832535 - INS CCTAATTAAAGATATTTCAACAGCAGAACAAGTAAAGTGGAAATGTTACATTGATTCTTCTTATGGTAGGAGATATTGGTTATATAAGACTGATCCTTTCCTGAATCGTGATGACTTGGATTCTAAGTCAAATTTAACGAGGTATGATTTGAGGGTCACAAAATCATAGAAATTATAAACCAGCCGGATTTCCTAAAGTTTGCCCAAAGTAAAATCATGCTTGGATGTGGTCTAGTTCCTCAAAGTGGTATTAGACGTAAACTATGTTACAGAGATTTAAAGCCACCAGTTTCTCAATTCTTAAATAGAAAAGGTGCGATCAGCCTTGGTGATACTCCACTACCAATAATTACCCCAACATTACCTCGTGGTGGGTGG tpg|BK006945.2|:831263-833305 7X173= 189=7X 
 tpg|BK006947.3| 300326 + tpg|BK006947.3| 300333 - INS ATATGTAATTATTTATTTACTTTTTCTGCCTCCTTGATATTAAAGTATTACACACTTTGACTTCTTTTTCTTCTTGTCGTTTCTCGTCTTTGGTTTAGCTTGCTTGTTGTGATGATTATTTGAGGCAATTTTACTACCTTTGCTTTTTGATTG tpg|BK006947.3|:300006-300653 7X5=71S 73S4=7X 
 tpg|BK006947.3| 583620 + tpg|BK006947.3| 583923 - INS GCCAACATTTCCAAAACGGATCATCACCACCATAATGATTGAATTTACAGGCTTAACGGTTTTTAAATTTATTCTTCGCATGATTAAATTGCAGATGCTGGTCTAAGATACAAAGTATGTAGCAGAAACTTTATCCATTGTTCGTGGTACTTGTCCCAATGATCGTATAATGTAATTTGCTCTTGAATCGTATCCATAACCTCCTCAAGATCTACAAGAGAT tpg|BK006947.3|:583162-584381 10S142=21S 52S4=7X 
 tpg|BK006945.2| 789512 + tpg|BK006945.2| 789621 - INS AAAGGAAATTCAAAATCTGTCTATTTATAGGCCGTCGCGCTCTACGAAAACGCGAAATTATTCAAACGGAAAACGGAAAAAAATCTAAAAAAAGAAATTAATTGAGAGATCTCACGGAAATGCCGCGAGGAATGTTTCTCGAGGCTGAGCGGCGTGGTCTGTGCAAAAAAATGGCAATTTTTTTGTAGGAGTTTGCATTGGGCCATTCAGAAGGAACACCGTTAGATGGGATGGTAAATGAATTTGCTGTTTCAGATTTGAATCAATCTTTACC tpg|BK006945.2|:788950-790183 7X137= 237S4=7X 
 tpg|BK006947.3| 688117 + tpg|BK006947.3| 688329 - INS AAGATGTTGTTCAGAATTTGTCATGTCATCTTCTGTGATTAGTGAAAATACGGGTGAATGGTCTATCATTGCTTTACCAAACTCCGCATCCCAGGTATTCACTCATTATGGAGCTATGAAAAAGACTACAGTTCATTATTGGCAAGATAGTGAAATTAGTTACACCTTGTTGAAAAAGTGTCTAGATGGTCAAGATTCGGATTTGCCTGGCTCCCTTGAGGTAATACAT tpg|BK006947.3|:687645-688801 7X47=1X166= 201=7X 
 tpg|BK006936.2| 726702 + tpg|BK006936.2| 726725 - INS TTTTTGTGTCGTTGGTATTTAGGGACGGTTGGTTACAGTGGCAATAATTGGAAAGTTCTTTCACAACAACACAAAAAAGGTGGAGAGAATAATTTGTACGGAAAAAGTTATACCTTTGCATGTCACGTGAACCAACAGAACATGGTAATACAT tpg|BK006936.2|:726382-727045 7X7=69S 71S6=7X 
 tpg|BK006947.3| 352984 + tpg|BK006947.3| 352694 - INS CTCTTCGTCATGTTTTTCTCTTCTGATACGCCTTTCCCTCCGCAGGAAATGAAAGATGAACCACCCATTACATTCGATTTTTTTTTTAATTATATTTTTGACTATTATTTAATCATTAAAAACACATATATTTCATAAATTCGTAAGGTCGTTAGTTCTATCGTAAAAGTGAAAAAGTTTTGAGCCAGTTTTCAAAAACCCGCAGGATCCCACTATGTATGGCTTTAAATAATGGTTTTTCACGTGCATCAAGTCCGTACTATCT tpg|BK006947.3|:352150-353528 7X4=145S 133=7X 
 tpg|BK006947.3| 333286 + tpg|BK006947.3| 333835 - INS GCAACAACAGCAATCCTCTGTTAAATACAGAGGATGTTACTAGATTTTACATGGCTGAGTGTATTTTGGCCATCGAAACCATTCATAAATTAGGATTCATTCACAGAGATATTAAACCAGATAATATTTTGATCGATATTAGAGGTCATATAAAATTATCTGATTTCGGGTTGTCTACGGG tpg|BK006947.3|:332910-334211 23S71= 3S156=7X 
 tpg|BK006936.2| 510307 + tpg|BK006936.2| 510634 - INS ATTGAAAATGGGGCTGACTTCGTGCCAAATCATTACATATTGTCAATGAGAAAGTCATTTGACCAATTGAAAATGAATGAACAAGCAGACGCTGACTTAGGAAAAACATTCTTCACTTTAGCCCAATTGGCGAGAAACAACGCTAGGCTAGATATAGCCTCCGAATCATTAATGCATTGTTTGGAAAGGCGGTTGCCTCAGGCAGAGTTGGAG tpg|BK006936.2|:509867-511074 7X14=63S 200=7X 
 tpg|BK006936.2| 675738 + tpg|BK006936.2| 676455 - INS CTATTACTCCTAACCATTTCCGTTTCTGATTGACCAGGCTCCGTGACAGGTTTGACTAATAGACCTGAATTACTCCAGTAAAATTGGTTATCGATATGATACAATTCAGCAAATTCAGGGTGTTCAATAAACATTGGATTCATTATCGGAAATCCAGTGACACTTGATTTATGAAACATGGTGTATAAGGTAGGTAGCAGGAAATATCTCAATTGGATAATAT tpg|BK006936.2|:675278-676915 7X7=104S 106S6=7X 
 tpg|BK006947.3| 263383 + tpg|BK006947.3| 263553 - INS ACAATGCATAAGGTCTTTTCCGGCTTCAAATATTCCAGCCAGTTTCCCTCATCTTGAGACAGGACAGGAACTTTGAAAAAATTCAATTGGTGAACCAGCTGTTTGTAGAATTCAGTGCGCTCGCTTCTCTTGGGGTAGAAAACAACAGGGTTGTAACC tpg|BK006947.3|:263053-263883 7X4=75S 74S5=7X 
 tpg|BK006936.2| 373199 + tpg|BK006936.2| 372752 - INS TTCTGTTGAAGGGTATAGTTATGCAATAGCAATTATTGTTACTGATTGAATGCCTTTATAATTTCGGTCCGAACAAAGTTAGGCAAGCGAGAATAATTGACGTTTGAAAGAGGGCTGCCAATGTACTATTTATATTAAATGGTGAATGAAGCAACGCAGTACCTC tpg|BK006936.2|:372408-373543 7X5=283S 145=7X 
 tpg|BK006947.3| 41158 + tpg|BK006947.3| 41409 - INS GTGGGGACGCAGATTGGAACTTGAAGACGCGATTTCAACCCACCAAGGGAAATCTATTAATGGCGATTTCAAAAGATAAATCGTGTCGTGTGTTCGACATTAGATACAGTATGAAGGAACTAATGTGTGTAAGAGATGAAACGGATTATATGACACTAGAATGGCACCCAATAAATGAATCTATGTTCACTCTGGCGTGCTATGAC tpg|BK006947.3|:40732-41835 7X4=182S 181=7X 
 tpg|BK006947.3| 192543 + tpg|BK006947.3| 192327 - INS TAAAATCTTTCAGTTTGTTTCAAAATGTATGTCCTTTTATCAGAATAAGTCAAAAGGGATGATGCCTCAAATAGCATCGGATACTAAAAGGACCGTACAACTTACCTCAAAAGCAGTGAAGTTGTCGCT tpg|BK006947.3|:192055-192815 7X112= 16S2=148S 
 tpg|BK006936.2| 392308 + tpg|BK006936.2| 392012 - INS GGACAGTATACCTCTCTCTCTCCATATTCACCTGTTACCCAGAGGGCACCATTCATATCATTATCAACGTAAAATCTGCGAATTACCGTAAACCGCAAAAAAAAAAGGATGGCGGGCAGTATCATCCTTCACGACCCGGGTGGCTGCTGCGCCCTCGCGAAAAAGAAATGAAATGGAGTGCAAAAACGGGAAAGACGCGCCACCGTTTCTGGCCCACGCGCTCATTCTCAGTGGCCAGGCACTAGAGACAGGACTGAAACCGCGTTACCACAACAAACAAAGGCAACGTGCAGTAAACAACC tpg|BK006936.2|:391394-392926 7X179=1D23= 284=7X 
 tpg|BK006947.3| 103229 + tpg|BK006947.3| 103283 - INS TGTTGGAATAAAAATCCACTATCGTCTATCCAAACAATTCTCTCAAAATTCGCCCAATTCTCAAAATTCACCCATTTCCCACACATATGTGTTTTAGGAACGTTTAGGATAAGGAATCGTCATACTGACGTACCTCATTTTGAGATACAACAAATCATATATTATAAGACTCCATGGCCAAGTTGGTTAAGGCGTGCGACTGTTAATCGCAAGATCGTGAGTTCA tpg|BK006947.3|:102765-103747 7X4=108S 105S8=7X 
 tpg|BK006936.2| 467419 + tpg|BK006936.2| 467649 - INS AACCCACACAGCACAAAATGTGTTACTCCTCGAAAAAATCTGTTACCCTTTTCCCGCCATGGTTGCCAGGGAAACAGTGGGGACTTCTGCGTTGCTTCTATTTTTCCCCCCTCCTTCCTCCTGCGCCTCCGTTTCTTTTTCTTCCCTTTTCATTTCCCTTT tpg|BK006936.2|:467083-467985 7X5=75S 76S5=7X 
 tpg|BK006947.3| 421686 + tpg|BK006947.3| 421905 - INS TATTTATATGCCAATGGATGCAGGTTTTCACCTTTATATATGATTCTATCAGTCCAAGACGGAGTTCTCGCCTTTTCAGAAGTATCATAATTATCTGTGCCATAATCATATTTATAGGTCGGACGGAATTGGAGGGTCGGTTCTTTAAAGCCCTGAAATACCACTCCTTCATTTATTTCTTGAGTCAACTGATCATATTGAAGCAATCTATCAATATAGCCA tpg|BK006947.3|:421228-422363 7X5=128S 111=7X 
 tpg|BK006947.3| 477657 + tpg|BK006947.3| 477624 - INS CCTTCAAATGAGAAACCCTGGTGTGTTCACGTAGATGCACAGACGGTGGGCAACCCAAAACTTAGTCTTCCGATAAACTTTTCAGGTTCTTGTACACGTGGAAACGCCCGATATATATCACATGTAGCTGTGTAATATGAGAATGCCTTTGTCCATGTGATAAACCGTGCAAAACTTAACATGGGAGCAGGCACAAGTGTGAGTCCCACGAACAAAACGCCGCTCGGGTAATAA tpg|BK006947.3|:477142-478139 12S21=91S 112S5=7X 
 tpg|BK006936.2| 611527 + tpg|BK006936.2| 611380 - INS GGGTTCTCATGCGAAATTATTTAAAGATGACCATTTTATATGACCCAACGTGGATATTTTGCTAATATATATGGTCTCATCTTCAGGTTTTTGGGAAGATGTAAATGAGGATAACAAGATGCGATGCTCATCCGAAGTGGTATCTAAATCAGGAAAGAACTGGCACGTTAAGGACGGCCACTTTGTTGAATTCGTGTTTAGGTAATCATAAAGTAGTTTAGTGTTTTTCTTCCAGTGCGAGTATCTTTCTTGCAAATCGATGGGTATACTGGAGGCTTCATGAGTTATGTCC tpg|BK006936.2|:610782-612125 7X518= 274=7X 
 tpg|BK006947.3| 402310 + tpg|BK006947.3| 402249 - INS GCCATAATGTGGGGACATTCCATGACAAAGCTATCTGAAGTAATTATTTCTCTTGTGGTAAAAGGTAAAGGTTCTCAAATAGCGACGTTTCTAGACTCGGAATCATTTGATACTTTGAATAATAAACCATGTAAGTATAAAAACCTATATCCTATGAAAGATCTATTA tpg|BK006947.3|:401899-402660 7X4=80S 79S5=7X 
 tpg|BK006945.2| 1035194 + tpg|BK006945.2| 1035000 - INS GGTTTGCAAGAACATGATTTGCTTTTTATGAGATTTCGGACAACTACCGGTGACGCAATGGGTATGAACATGATATCGAAAGGTGTCGAATACTCTTTGAAACAAATGGTAGAAGAATATGGTTGGGAAGATATGGAAGTTGTCTCCGTATCTGGTAACTATTGTACTGATA tpg|BK006945.2|:1034642-1035552 7X281= 151=7X 
 tpg|BK006947.3| 407773 + tpg|BK006947.3| 407191 - INS TGTACACATTCTAGTGGGTTGAATTGCGGACGTTGGGACTATATTTTCTCTACAATCAAGAGATTAAGAAATGATCCTAATCACATTTTGCCCAATAGAAATCAAGTGACTATGACTTCCCCATTCATGGATGCATACGTGAAAAGATTAATCAATACCTGTCATCGGAGGGGTGTTCATGCC tpg|BK006947.3|:406811-408153 7X3=103S 92=7X 
 tpg|BK006947.3| 376055 + tpg|BK006947.3| 376341 - INS CAAGAATCCCGTCACTGATCAGGAATGGTGTTCAAACCAAACAAAGGTCCATATTTGTCATCGTTGGGGACAGGGCACGTAACCAGCTCCCAAATTTACATTATTTGATGATGAGTGCTGACCTTAAGATGAACAAGTCCGTCTTATGGGCTTATAAGAAGAAGCTTCTAGGATTCACTTCGCACAGAAAAAAAAGAGAG tpg|BK006947.3|:375641-376755 7X7=93S 92S8=7X 
 tpg|BK006936.2| 756271 + tpg|BK006936.2| 756807 - INS CTTATAAGGTTGTTGCGTATAATACCGTCTATATTCTGGAAGACTTTGCATTAGCCTGCTTCCTGTATCTTCTGGATATAAATTCTTGTTAATAGCTGATAAATCAAATTGTTTATTCTCGCAATCACTTGAAGACGCTAGCTTTCGCCTCTTTGGCGTTGGCGATAGATCGCTTTGTATATGCATATGAGCTTGTGGAGATGGAGGTGGCAAGTTAGTTTTCATCCACGGAGAGCTTCCATTGGAATAATTATCGTGTTGAGACCTACGGAGGATATGC tpg|BK006936.2|:755697-757381 7X87= 13S246=7X 
 tpg|BK006947.3| 29705 + tpg|BK006947.3| 30346 - INS GCTTTAGCAACATGACCTTTATTGTTAACACCACGCTTTAGAAAGCGTGCACCAGCAAAATGGTGGGATCTTCTTGCGATTAAAGTAATATATATGGACTTACCCAAAACTGAAACATTAACCTGGTCAATAAATCCATGTATAATGCATTGGAAC tpg|BK006947.3|:29379-30672 7X1=2I75= 154S4=7X 
 tpg|BK006936.2| 274642 + tpg|BK006936.2| 274974 - INS ATTCTATTCTTGTCAATAAAGTGGAAATGTGTCAGATGTCACAGTTTCTTTATTTGTGACACATATTTTCAACATAAATTCAGGCATTAGTGCTTTTATAAGCATAAGAAGTTGTGGCGATATGAATATTCCAGATTTTACTTACAAGCTGCATTGTATTCCTAAAATTCTTTTTTCTTTTTTTTTTTTTTTATG tpg|BK006936.2|:274238-275378 7X6=91S 24S12=69S 
 tpg|BK006945.2| 265565 + tpg|BK006945.2| 266068 - INS ATAGAAGATAGTTTACATATCAAATCAAAAAAATATGATATCAAATTTGTATTGTCGTTCAAGTCTATACCTTGTTTTACTACGCGATTGCCATCATATTTGGGCTTACCGGATAGCACAATGATATACAGAGCAACGAACATAGGAACGTTCAAAGCCACCAGCTTAATCCATTGGCCAATTGTAACCT tpg|BK006945.2|:265171-266462 7X9=86S 89S6=7X 
 tpg|BK006947.3| 492792 + tpg|BK006947.3| 493162 - INS CTCCAAACTTTTGAAATTGAGACAGTCCTTGAACGCTACAGCAAACGACAAGTACAAACTGTCCATTAATGACCTATTAGTAAAAGCCATCACTGTTGCGGCTAAGAGGGTGCCAGATGCCAATGCCTACTGGTTACCTAATGAGAACGTTATCCGTAAATTCAAGAATGTCGATGTCTCAGTCGCTGTTGCCACACCAA tpg|BK006947.3|:492378-493576 7X2=160S 100=7X 
 tpg|BK006947.3| 162105 + tpg|BK006947.3| 162164 - INS AAACTTGAGATTCTTTTTCCATCTGTTCAAACTTTACTAAAATCTCTTCGTTACTATTTGGGTTTTTTATAGCCTTGTTTTCTAACAGATATTGCAACTTAGATGCAATAAGCTTATAGTC tpg|BK006947.3|:161849-162420 7X4=20S 61=7X 
 tpg|BK006936.2| 84444 + tpg|BK006936.2| 85005 - INS AAATAGAACATCAATTAGCGTCGATATCAAAGGTAACATCAATTTGAGGCACACCTCTGGGAGCAGGCGGAATGCCACTTAATTCGAATTTACCAAGTAAGTTATTATCCTTTGTTCTTGTTCTTTCACCTTCAAAGACTTGAATTAAAACACCAGGTTGATTATCTGCATAGGTAG tpg|BK006936.2|:84076-85373 7X4=251S 155=7X 
 tpg|BK006947.3| 513617 + tpg|BK006947.3| 514366 - INS GCTTCCACAACTGATGACCAAACCTGTTTTATTTCCGCTTGGGTTATAATTGTAAAAACTAAACAGACTGTCTATTCCGAAAGTAACGCCTGGTACATTGTAAGTTTCAAACAAAATCTGGTACCAATTTGTCCGTTGTGATTGAACAGTTGCCAGTCTTTCGGTAAGTAATATTGGATTAGGAATTCCGTTATCTGGTACCACTCCCAAATGATGAAAAGTGTAGTCCAATATTTCTTCAGTGAGATTCCAATTGGTTACAAATGGTCCGTCAAAGGGGCTTCTCGATTGCGAACGCACAGCT tpg|BK006947.3|:512995-514988 7X116= 152=7X 
 tpg|BK006945.2| 565637 + tpg|BK006945.2| 566066 - INS CCTTGTCGATCTATCTAAGAGGTTGTCGGAATCCATCATAATAGCCCTTGGCGTAAACTTATTCCTACTGTTTTCGCGGAAGAAAGGCTTTGTGTCATCATCTCTTTCCGTACTGGAATCAGGAAGCTGAGATAGCCCATCGGTGCCTATAGCGTGTTCTTTCGCCAATTGAGACCAGAGAAACTTACCAACGTGGTTCCCGCATTGACCTGCTTGCAAAGTAATAATTTCTCCACCCATAGATAGTTATATGTTGAATTCTTATACATGTGACTAACCGATATTACGCATTTGTTCATTTCGCAGCTACTGTTACGATTATTATTTATTACATTTAATGAAATTTCCCAAAAGATAATATTAACGCGTTCTGTTACCC tpg|BK006945.2|:564865-566838 7X12=184S 2S354=7X 
 tpg|BK006936.2| 81725 + tpg|BK006936.2| 82069 - INS TTTCTTTGAAACAACCTCCTTAACACCCTCTTCTTTGAATTTCAAACTTTCAGCTTTTAAAACAGGTGAGTTTATCAAGTACAATCTTAATGCATCCGCACCATATTTGTTCAGAACAATGGATGGATCAGGGTAATTTTTCAAGGATTTAGACATCTTTCTACCATCGGCAGCTAAGACAATACCAGAGACGATGACGGTCTTGTATGGAACAGAGCCAAATAGATGGGTACCTAAGACAGCTAACGTGTAGAACCAACCTCTTGTTTGATCCAAACCTTCAGAGATGAAATTAGCTGGAACTCTTTCGTCAAATTTTTCTGTGTTTTCAAATGGATAATGTTGAGAAGCATAAGGCATAGAACCAGATTC tpg|BK006936.2|:80967-82827 7X288= 13=1X172=7X 
 tpg|BK006947.3| 35838 + tpg|BK006947.3| 36236 - INS ACAACCCTGCTAGCGCTGGTGTCTCTTCCGCATTGTTAATATTTTCCATGATTGTAATGTTTGTCCCCACCGTTTTATACGAGATATATGGCGGCTACTCGGTAAACTGTGCAGACGGTGCTAACGACCGTGACTGTACTTTCTCGCATCCTCCCCTGAAGTTCAACCGTTTATTCACTCATGTTATTCAACCTATGTCCATATCTTGTGCCATTGTTCTCTTCTGTGCTTATATCATTGGCTTGTGGTTCACCCTTAGAAC tpg|BK006947.3|:35300-36774 7X215=22S 1S1=25S 
 tpg|BK006947.3| 579038 + tpg|BK006947.3| 578794 - INS CTGTAACATATCC tpg|BK006947.3|:578754-579078 7X3=3S 7=7X 
 tpg|BK006947.3| 17137 + tpg|BK006947.3| 17385 - INS TAGTTGGCACATGTAAACTACG tpg|BK006947.3|:17079-17443 7X5=6S 7S4=7X 
 tpg|BK006947.3| 511554 + tpg|BK006947.3| 511414 - INS GCTAATATCAGCTATGATGAAAAACACAGGTTGTGTTTTCGCTAACGACGCCAATAAATCTAGAACAAAATCTTTAATTGCTAATATCCACCGTCTAGGCTGTACCAACACTATTGTATGCAATTACGATGCCCGTGAGTTCCCTAAGGTAATTGGAGGTTTTGACAGAATTTTACTGGATGCCCCATGTTCCGGTACTGGTGTTATCGGTAAGGATCAATCTGTCAAGGTGTCTCGTAC tpg|BK006947.3|:510920-512048 42S248= 120=7X 
 tpg|BK006947.3| 325151 + tpg|BK006947.3| 325623 - INS ATGGCATCCTACATGAACCAACAAACTATTGAAGAGTTTGATTCTTACAGCCGTTCCCGTCCCACAAGACCGCTGGGTTATCTCCCAGTATGGGCCAGATACACAGATGATAAAGTTAGTGTCATACCGAAAAAAAGAACTTTGAGAGTAGCTACCTTGTACTTACAAGAAACTGATTCGTTTGATGATGGCTCTAGTTTAACATCTACCAATTATACTGAAATGGGCTCTAATATC tpg|BK006947.3|:324663-326111 7X2=164S 119=7X 
 tpg|BK006947.3| 612391 + tpg|BK006947.3| 612892 - INS GTGCTATGCTATTTCATTCCATTCTTTCTTAGCTAATAACTTATCATTAGGTAGCCTATGGCCAAACAACTCGACAAGCTGTTCATCTTGAAGTAGTCTCACTATTCTAGATCTGATATCACCAATTGCTGGGCCACCAACTATTCGTAGAATTTCACTTGTGGACCCGCCATTATCTGATATTGGCAATATATACGTCAGCTCATGTCCTTTTAAGATAGAAATATTAGAAAAGCAAGGAGTCAATGAATTTGTGGCAGTCCCACCGGAGCACACAACGACGTTCATCTAGTAAACTATCTCACCACACTCTGCTATTTTGTCCCCTTATTACCTCGAGGGAACAAAAGATTCCGTTTCCTCTCTTTCATAGTCCGCCTAAAT tpg|BK006947.3|:611609-613674 7X5=172S 360=7X 
 tpg|BK006947.3| 526333 + tpg|BK006947.3| 526165 - INS TAGAGAAGAAGAAACCTGCCGTCATCTCCAATAATATGCCTACAAGTAACATTGCCCTTTATCAAACAGCGAGATCGGCGAATATTCATGGTCCATCATCAACTTCCGCATCTAAAGCGTTCAGAAAGGCTTCGGCCTTCTCCAATAACACGGCACCCAGCACTAGTA tpg|BK006947.3|:525815-526683 11S92=30S 37S5=7X 
 tpg|BK006945.2| 387419 + tpg|BK006945.2| 387607 - INS TCCGTACCAAAAGGAGAAGAATATGTGTTTGATCTAAATGTAGAAGAGCCCGAAGTGGAAAATGTCCCGTATTGTTGACAGTCCATGTTTGCTTCCGAAGCAGGCACGGATTGAGTTGCCGTACCTGAACCGCCTCCTAAGCCCGTAGCAGTGGGGCCAATGGCACTGCCCGTTCCCGTCAACCAGCCAAATGGGTTTATATCATTAATCAAAGATCCGCCGCTTGACGAATCATCACGTTTGTCAATAACACGTCTCCGGCTACTACCCATAC tpg|BK006945.2|:386857-388169 7X171= 8S62=1X1=1X184=7X 
 tpg|BK006947.3| 424845 + tpg|BK006947.3| 425268 - INS GTCCTCTTCTCTACATCCTTCTACACGGTCGGCACCTGCAAGCATACCTAACTCTGTGGCGGCGACACCGCAACCACGGTCATTGTGACAATGTGTAGAGATGCAAACCTTCTCACGCTCAGTAATATGGGTAGCGAAGTATTCAATCTGATCAGCATAAACA tpg|BK006947.3|:424505-425608 7X5=76S 77S5=7X 
 tpg|BK006947.3| 285305 + tpg|BK006947.3| 285582 - INS TTGATGTCGTCATTCAAGCCGGTGTTGTTCCAAGATTAGTAGAATTTATGCGTGAAAACCAACCTGAAATGTTACAATTGGAGGCTGCTTGGGCTTTGACTAACATTGCATCAGGTACATCTGCTCAAACAAAAGTGGTTGTTGATGCTGACGCTGTA tpg|BK006947.3|:284975-285912 7X6=73S 73S6=7X 
 tpg|BK006945.2| 196979 + tpg|BK006945.2| 197049 - INS TCTCTAAAGTTTTTGTTTCTTTTCTTGTAACTCAACACACTTTGTTGAAATTCTGAAGTTCTATCCTTTATGTTCATGGGAGTTGTGTGGTATGGTGAAATGGTCGTTGGAAACAGAGGTGGAATAAAATATATACAGTAAAGAGTGGGTGATTTCCGTTCAAAGGTCTAACAGGAGCGTCGATGCGGCGGTAGGATTTTTTTTTTTTTTTCAATTTCTATATTGACATTATTATCATAATGATTGTTTCGAATATGCCCTTTCGCCTCGCCTCGATCAATAAACCT tpg|BK006945.2|:196391-197637 7X6=466S 144=7X 
 tpg|BK006947.3| 499612 + tpg|BK006947.3| 499778 - INS GTGTCAACAACGTCCCAGTTAGAGATGGTGTTACTATCGAATTCTCTACTAACGTAAAGGACGAAATCGTCTTATCTGGTAACTCTGTTGAAGACGTTTCCCAAAATGCCGCTGACTTGCAACAAATCTGTCGTGTTAGAAACAAGGATATCCGTAAGTTTTTGGATGGTATCTACG tpg|BK006947.3|:499244-500146 15S80= 14=82S 
 tpg|BK006947.3| 44202 + tpg|BK006947.3| 43717 - INS CAACTGCAACTGCACTCAGATTGAACTTGTCTAGGAAGTGGCAACACGAATATAGGGTTATTCCTGGCATTTGCCATCATCTTATCATAAACGGAGACAGGAATCACAGCGCATAATGTATTATCTTTTTGTGCCCATCTTGCTCTCCAAAGAAACTCTACTTCCTGTTTCGATAAGTCCTTCAG tpg|BK006947.3|:43333-44586 7X5=216S 3S171=7X 
 tpg|BK006947.3| 615420 + tpg|BK006947.3| 615062 - INS GAATTTAATGACGTCCATATTGATTACACCTGATGGTAAAACGTTTGAAAGCGAGGCTGCCCATGGTACGGTGACCAGACATTTTAGAAAACATCAAAGAGGCGAAGAAACATCAACAAATTCAATAGCCTCAATATTTGCCTGGACAAGGGC tpg|BK006947.3|:614742-615740 7X1=2I54=19S 7S1=152S 
 tpg|BK006947.3| 397329 + tpg|BK006947.3| 397074 - INS TCTGTAAGTATTCCAAGTAATTTAATTCCGAGGTACCGTGCCACTAATTTAGAAGCTATATCTATCGACTGCAACGTTAGCACCAGATGTAATTCCGGTATTTTGACAGATAATGATGGTACAG tpg|BK006947.3|:396812-397591 7X5=57S 50S12=7X 
 tpg|BK006947.3| 10026 + tpg|BK006947.3| 10661 - INS GATGTATACTGATCTTAATCACGGATGTATACTGATAATAGGGTTGACTGCGCCTGTACGGATTACAGTGCCCTCTTCAATTGGAAAATCCAAGCTTTCAAGATGCGTAACTGTTATTCAAAGGATCCTCTAAGATAAAACACAGATCGGCAGATCCGAGAGTTGGCTTCTGTGCCTTGGGCTCAAATTCCTTTCCCACCTCATTCAAATTGATTTTTCTGACTCCAAAAAAAGACAAAGCCCTGCGATAGTTCCCGAATGTTGTAACATCAAAGC tpg|BK006947.3|:9460-11227 7X8=2S 259=7X 
 tpg|BK006947.3| 227631 + tpg|BK006947.3| 227672 - INS ACGTATAGGAGTGATATACATGCAGAGGTGGCTACAACTGTGGAAAATGGATTTGGTACAAAAAGTGTCTCATGGCGTTTTTGAAGGCTCGTCCGAAGAACCGGCTGCTCTTATGAATCATGATTATATAGTAT tpg|BK006947.3|:227349-227954 7X3=16S 67=7X 
 tpg|BK006947.3| 399015 + tpg|BK006947.3| 399033 - INS ATACTGGAACATGCAAAATCGTTCTTG tpg|BK006947.3|:398947-399101 7X4=9S 8S6=7X 
 tpg|BK006945.2| 637241 + tpg|BK006945.2| 637422 - INS TTTCTACTACTTTGCAAGTCGTTAACGAATTGTTGAAGGACGAAACCGTTGCTCCAAGATTTAAGATTGTCGTCGAGTACATTGCCGCCATTGGTGCTGATTTGATCGATGAAAGAATCATTGACCAACAAGCTTGGTTCACCCACATCACCCCATACATGAC tpg|BK006945.2|:636901-637762 7X5=76S 76S6=7X 
 tpg|BK006945.2| 180998 + tpg|BK006945.2| 181646 - INS TTATTGCCACTGTCATCATCATTCTTGGCAATAGGAAACCATGTCTTTTTATCTGGAAAAATTTTCTCTGCACCCTTCTTAAAACTTAGCTTATTAGGAAGAGGTGACAACCACCATTGCATTAGTTTGACGGAAATATGGACTGGTGAAAATAAGAAATTTCGGTCCCTTAAAACTCTATCCCATAAGAC tpg|BK006945.2|:180602-182042 7X5=90S 91S5=7X 
 tpg|BK006945.2| 779273 + tpg|BK006945.2| 779807 - INS CTCCAATGATAACCTGGCTACTTTTACCACCGAGAAGCTTGATGCTGATGGTGGGCATGTTCCTTTTAACGTATCACTCACCATGGTCTAAAGTAGCAAGAAGGCTTTTATGGAAGTTTAAGATTGTCAGGCTGCTTGTTTTCTACGTCACGGGTTTAGACCTTGGTGGAATAAATAAGGACCAGGGTATTTTTGCTACAGTGCAGAAGCAAGTGAAAAAGTTGGCATCAACAGAAAACAGTAATGGCGTATTATCCGATTCCAAGCC tpg|BK006945.2|:778723-780357 7X131=1X32= 134=7X 
 tpg|BK006945.2| 985802 + tpg|BK006945.2| 985996 - INS ATTCTGAATAAGGTGAGATTCTTCAAAATTGCTGATGATTTTGGTAACTCAAAACATTTATTTTTTGAAAGAAAGGGGAAGATAGTTATATTAACACCAGAATTTGATCAATTGACAAACCAAGTAAAATATTTCAAATTTTACAAAGAGTATAAGCTCCCAAGTTCAAGTAATAACATTCTGAATAACGAAATTGAGGATATTGCCATATTCAGGAAAAGTTTTGCTGTGTGTACAAAGAAAACAGTCATACTTTATCAAGATTCATTCGAGGATAACGGAATAGTCTTACCATCTTTTTTGAATGATAAAGATATGATGGCACACTTGAGGCATCCACATTTGAATAGCTTACCGTTCAAAAGTGCTACAGACTCCAAGAAACGCCCCTCCATAGAATCTCTCACTGAAGAAGCAAAAAAGGATATCGCCACTTGCAAAGCTATAC tpg|BK006945.2|:984892-986906 7X260= 224=7X 
 tpg|BK006936.2| 241339 + tpg|BK006936.2| 240600 - INS TCCTATCTATATGTTCCCCTAACATTTACATGTTTGAAACCGTTGGAATTGGCCGTCCCGACTTTAATAACTTTGGGCCCAGTGTCTTCTATGGTAATTTGGTGATTCTTGTCTGTGTCCTCACTAGCGAGCAGCTCATCTAAAGCGAGATCCACATTATCAATATAAAATCTACGGTTACCTTGGCTGCTGAGGAAGCTGTCGTCTTCAGAAC tpg|BK006936.2|:240158-241781 7X6=147S 107=7X 
 tpg|BK006936.2| 425335 + tpg|BK006936.2| 425308 - INS GTGGAAACCCTGAATACCACGAATAAATCGTCCATAATTGAATACTCAAGTGTTTTTGACGAAAGATTATCACTTGGAAACAAAGCAATATTCCATTTGGAAGGGTTCATAGCAAAAGTTATGTGCTGTCTAGATTAATGTAAGATATGTCATAAAT tpg|BK006936.2|:424980-425663 7X5=73S 73S6=7X 
 tpg|BK006936.2| 797513 + tpg|BK006936.2| 797925 - INS TCTGTAGAAGAAACTGGCATTCCGATTGCAGTAGCAAATGTTAACCAACAAGACGAGCCAATCAAAGCACTGGTCATAGTAAGCATTAAAACAGCGGGGTCGTTGGTAAAAATGGAGGAATCTATAATGTTGTTCTTGATAGTACCAGAAACTCTTGCGCCTGCCAAGACAGCACC tpg|BK006936.2|:797147-798291 7X1=1X5=1X108=16S 1S1=434S 
 tpg|BK006936.2| 536078 + tpg|BK006936.2| 536276 - INS GCCCAGAAGGATCGTCCCAAAGCTAGCCACATTTTATTCGGCGAATCCTAA tpg|BK006936.2|:535962-536392 7X6=19S 23S3=7X 
 tpg|BK006936.2| 738392 + tpg|BK006936.2| 738461 - INS ACTGGAAGGAGGAATTCGCCAAAAAATATGATAATGAGGCTGAAAACACAAAGATTATTATCGTCAGTAGGTCAGAGGCTAGACTGCTGGACACATGCAACGAAATTAGGATTGAAGCTCACCTGAGAAGGGAAACCACTGACGAGGGCCAAGTGCAACATAAGTTGGCTGCGCCCTTGGACCTTGAGCAACGGTTATTTTACTACCCATGCGACTTGTCCTGCTACGAATCCGTGGAATGTTTGTTCAATGCCCTGAGAGACTTGGATTT tpg|BK006936.2|:737836-739017 20S182= 13=1X241=7X 
 tpg|BK006936.2| 111691 + tpg|BK006936.2| 112365 - INS AGAGGAAGCACAGATTAAAGCTCTTAATATATAAATGCACGTATATCTATACCCGTAGTATATATCATTTGTACCTCAATACAATTTCAAATCACCTGTTATTTGATCCAATACTGCTTTTGGAGCAGGTCCTAAACCCAATACGGTGGCACTTCCCGCAGCAATCTGTGTTCTACCAGCATCATGAATAACTGCTGCATTCACCCCAAGTGATATAG tpg|BK006936.2|:111241-112815 29S68=19S 105S4=7X 
 tpg|BK006936.2| 534382 + tpg|BK006936.2| 535157 - INS TCATGGAGTAGAAATTGGCTCGACATATTTAAAAATGTCGACGGGAAACTGAAACCAGGAGGAGTAGAAATTGGTTAAATTGATTAGCTAAAATTTACTCGTTGTGGACAGAGTTTGAGCCAAGCGGAATGTTTTCAAGGCTTTCTTTGTTTCGAAGGGCAGCTCTGGCTCCTGCCCCTATGAGAATGTCTTTTAGGACTATTTATCAAAAAACCGAGGATGAATTGCCCAGAAGGATCGTCCCAAAGCTAGCCACATT tpg|BK006936.2|:533850-535689 7X3=211S 10S6=1X9=1X216=7X 
 tpg|BK006936.2| 617938 + tpg|BK006936.2| 617794 - INS AATTCATAGCTCTAGGACAATTCTATTCAAGTCTGACGCCGAAAACGGACCATTGGACCTCCCCTGCTGTTGAGACTGGCCTTGACTCTGTTGCTGTGGCTGCTGGCCGGAATTGGCGCCAGCAGCATTATTAGTTCGTTGATTCTTTACTGGTTGTGGCTGATGCGTGCCATTTTGATTCTGATTCGTACTTTGCTTCTGTGACATTCTTATTTTTCAAGTATCTCAACTTGAACCCGGAG tpg|BK006936.2|:617296-618436 16S111=1S 116S5=7X 
 tpg|BK006936.2| 511629 + tpg|BK006936.2| 511833 - INS AAAGTCTACATGATAGGTGGCAGCACACCGCAGTAGATGGAAAACTCGAGTTTTACATGGAACAGGTAGATAAATTTCCTCCAATCTTGTACCAATGGTTTTTAGAAAACTTTCCTGATCCAATCAATTGGTTCAACGCCAGGAATACGTATGCC tpg|BK006936.2|:511305-512157 7X24=53S 3S1=200S 
 tpg|BK006945.2| 14287 + tpg|BK006945.2| 14204 - INS TATGTGTAGCATAATTTGTCCATTCTTTATCCGCATTCAGGCACTCCCAATCTTTATCTCTAAGGCAAAGAGCAACCACCATTTCACCTCTGGAGGATCTAGGCATAAAATATATTAGGCTCTCAAGGGAAATGAAGCGCGGCCGTCGTACACTCTTGGGCTTCCCAAGCCCTAGATTGAAATCAACGTCATACAGGCTGACTTTTGCCCACGAAC tpg|BK006945.2|:13758-14733 7X78=30S 6S1=318S 
 tpg|BK006945.2| 957002 + tpg|BK006945.2| 957299 - INS AATATTCATCCAACAATGAACAAATATTCGTAACTGTACCAATGAACCATCAATCTCAATTTCCGTTTCTTCATTCAATGGAAAACTATCTTGGGTACTACCATCACTGGATAGAGTTTCTACCATGGTTGCTTTCGTAATATCATCAGTAGACTGTCCCTCATTATTTTTTAGAACCAGTTTATCGC tpg|BK006945.2|:956612-957689 7X7=87S 90S4=7X 
 tpg|BK006945.2| 746657 + tpg|BK006945.2| 747105 - INS CAATTGACAATTTTGATGCTATTGTTTTTATAGTGTAATTGCTATGAGTTTATTTTGTTGACAAGTATACTTGGCTGTCTTTTTTATATAATAACGAAAATGTGTAGTGGAAAAGCAGGTGTGTTTTGTCTTATATCTTACAAACTATATAGGCTTATATAGTTTTTTTTCAAAGATTCTTATTACTGCACAAAAAAAAATAAGATCCCAAATTGAACATTAACATTAGTCATATTCAGGGATGGCTCATCACGAACAGCAAACTGAATAATTTTCTTGTCTGCGTTCCTTTTTTTGTGCACCAATGGATGTAGTATGCGCACCTGATGCGCATAATAGATTGCAATTACACTGACTACAACTTACG tpg|BK006945.2|:745909-747853 7X213= 184=7X 
 tpg|BK006945.2| 124103 + tpg|BK006945.2| 124388 - INS GTATAGGATTTGGAGTAGGGTAGTAAATATAAGGATTCTCCTGTTGCTGTTGCTGTTGTTGGTCTTCTTGTTGTTGTTGTTGTTGCTGTTGCTGTTGTTGCTGGGGAGCAGAGAGTGGTGGAGGTGGCATAAACATCATTGGGTTGGGGTAGGCAAACGGGAACGGAGAATTGTTTGGAGGGGACGAAGGTGAAGAAACAGAAGAAGGTCTGTTTGCCTTCTTCTTTTTCTTACCATTTGAGTCTTCGGTGTCTTCATTTGCTGGAATCTGTACTGAAATCATCTGGGAGATGAAATTTGAAGGAGATCCGATCAAGTAGTTGGGGAAGTTT tpg|BK006945.2|:123425-125066 7X3=195S 166=7X 
 tpg|BK006936.2| 639197 + tpg|BK006936.2| 639625 - INS AGTCTAACCCTGTAAAGAACAATCACGTTCGCCCAAAGCAATGGCCTTACCAAAACCATCTCCCATAAGTTGGACTTCAACATGCCTGGCATTTTCGATAAACCGTTCCAGAAATACACCAGCGTCACCGAAAAATGTTTCACCTTGATGTTTCACAGTCTCAAAAATATGCTCGATGTCCTCTTCAGAATCGACTTTCTGC tpg|BK006936.2|:638779-640043 98S100= 177=7X 
 tpg|BK006936.2| 497344 + tpg|BK006936.2| 498041 - INS GTCTATGGGAACGGAAGAGACGAAGAGGAATCACAGGAGCAACAGCGACGGGAGCACCAAGAGACTACGCAAAACAATACAAGCGAACTCTCTCTATCGGAAAGAGTGATACACAACGTAACACTCCCCATTTCTTTTGCATACGACGCTATACATGAAGTGAGTACCACGACTGGTGTTTCGGGTAGCTTATCCATGATAATGGACTATGTACCGAAGCCCCATTGGCCGTTCATTTCATCCTCTAACAAAAGTGCCGACAAAAATAATTACTCAAATAGCAATGATAACGCAAATTCGAATGCCCCACTGA tpg|BK006936.2|:496704-498681 7X186= 294=7X 
 tpg|BK006936.2| 40749 + tpg|BK006936.2| 40919 - INS AAACAGGTAAGTTATTGAGCGGGTTGGCACAAAGAAAGACGAATGGGGCATCTAACGGAGATGACAGTAACGGGGGAAATGGTGAAGGGCTTGGAGGTGACAGTGACGAAGCAAATATAGAGATTGATCCCTTAACTGGTATGCCTATATCTAATGATCCTGATG tpg|BK006936.2|:40405-41263 7X147=7S 1=165S 
 tpg|BK006936.2| 128031 + tpg|BK006936.2| 127265 - INS GTATAAGGAAGGGTAAATAGCACCTCTCTTCTTTTAGTGCTTTTTAGCGTATGATTCTTTTTAAGAATCTGGTCTTTCTTCCTTCTATTTTGATTGGGTATATTTCTATTCGTGTTTCATTACTGGTCTGGGTTAATTGGGTTTTGGTTTGGTCCAGTTGTTTTCAAGTAGCCTTTATTTTTTCATTGTGGTATTTTATCTTATCGATTTATACTTTTTTTTATTCAAAGAAAATTAAACAGATAATCTCTTATGAGCCTAGCTACTTTGTTTTTTCTTACAGGGCCATTGACT tpg|BK006936.2|:126663-128633 7X4=190S 10=1X265=7X 
 tpg|BK006936.2| 463969 + tpg|BK006936.2| 464433 - INS GTTCCATAGCTTGTGCCTTTAGAAGATAATCCAATGCCTTTTGAGGGTCATAAAATTGTACGTTACTCATACCGTAAAGACAACCTAATTGTTGTAATACTTTGGCATGATGTTGATTTTGAGCCAAGACATGCTCGTAGGCTTCCTTCGCACCTTGCCACTCTCCCATACTCTCCAAAACACTACCCAACTGAAACCATATGTC tpg|BK006936.2|:463545-464857 7X15=87S 99S4=7X 
 tpg|BK006945.2| 840729 + tpg|BK006945.2| 840029 - INS CCTCTTCTCTGGTCTTGGAGTTCACCACGTAATGCCTGTTTAAGACCATCAGTTAACTCTAGTATTATTTGGTCTTGGCTACTGGCCGTTTGCTATTATTCAAGTCTTTTGTGCCTTCCCGTCGGGTAAGGGAGTTATTTAGGGATACAGAATCTAACGAAAACTAAATCTCAATGATTAACTCCATTTAATCCTTTTTTGAAAGGCAAAAGAGGTCCCTTGTTCACTTACAACGTTCTTAGCCAAATTCGCTTATCACTTACTACTTCACGATATACAGAAGTAAAAACATATAAAAAGATGTCTGTTTGTTTAGCCATCACAAAAGGTATCGCAGTTTCTTCTATAGGCCTCTACTCTGGTCTTTTGGCTTCCGCTTCATTGATTACATCTACTACTCCACTAGAGGTTTTAACAGGATCCCTTACTCCCACTTTAACCACTTTGAAAAATGCGGCCACCGCCTTGGGAGCGTTTGCGTCAACTTTCTTTTGTGTGAGCTTTTTCGGCGCTCCTCCCTCATTGAG tpg|BK006945.2|:838961-841797 7X4=401S 511=7X 
 tpg|BK006936.2| 368585 + tpg|BK006936.2| 368684 - INS TTATACCCAATAATTGCGAAACTGTATCAGTTATTTTCCATTCAGGGATCGAGGCATCAATATTATACAGAAAAAATGATTTGGTGGAGGGGTTTTTTAAAAACGATTCATTCAAGGGTAGTTTCTTCAAAATATGAGAAATGTCCACGGACGCGTACTTTTCCAAGTTTTTGACCTCATTTGCACCTTTTTCATTTTTATACAATGCAGTTGTGTTTTTTATTAACGGAGTACTTGGGC tpg|BK006936.2|:368091-369178 7X188=22S 1S1=161S 
 tpg|BK006936.2| 708302 + tpg|BK006936.2| 708279 - INS GTGGTGTAGGATACAGGTGTCCTGCTTCTGAAGTAAAAGTCTAATTCGAATAGGGGACAATCTCTAATTTCATCACGCACTAATTCGTATACGTCATCTCTATCCAAGCCATACTTGAATAACATGAGAAGGATAAAACGATCTTCTTCTTCAGAGTACGTCCTTTTGTGGTTAGAAGAAGGAGGATGTTTTAATTTCAAATCGAAGAATGGATTCTTATACTCAGACAACTTCCGACGTAAAGCCTCTTGTTGCATTTTGACACGCTTGATCTTCTCTTCTTCATTCTCAATTATTTTCAGATATTTCTCATAATCTTCAATTCTTTCAATGTTAGACCAGAAGGCCTTAGCATATGCGCGAACTTCCTCTAGTGTTTTGCCAGGGGCCAATTCTCTCGCAATGGCTTGAATGGAGTTCCTACCGTATTTACCAG tpg|BK006936.2|:707393-709188 7X158=9S 156=1X266=7X 
 tpg|BK006936.2| 649172 + tpg|BK006936.2| 649070 - INS CTATAATACTCGCTCCATCCGACGGGCAACCAATTCTCCAATGCTACTAATAACTTACCTCAATTTGGGAACGCGATGTCAATTTCTATGCAACTGCCCAATGGCAACAGCAATAAAACGGCCTCAAGCATGAACACAAACCCTAACACAAACATGATCATGAATTCTAACATGAACATGAACATGAACGTAAATCCAGTACCATACGGAATGGGAAACGGTGCAAATATGTATGACGTGTCCAGGATGATGAC tpg|BK006936.2|:648548-649694 12S148=37S 57S7=7X 
 tpg|BK006936.2| 214436 + tpg|BK006936.2| 214722 - INS GGTAGTTCTCTGGCTCTTTTTCCACATACGCTAAATCTTCATTGGATAGTTTATCAGCGGCGACAGCAATCTTGACACCATTAGCCTTGTGCAAGTGGATTTTCCCCTTAGCACATCCAATGAATTCTGCATCCACTTTGAAAGTACCACTTCTATCAACCCATAGACGCGATTTTTTTGGATTGGGGAAATCTTTGGTCGCCGAAGAGTTTTTTTTGTGAGAGGACAATGAACTTTTTCTTGACCTTTTACCGGCAGCACTACCTACAACATCGTTTTGTAGTTCATCATCTTTCCAACTGGCATTGGCATTGGATTTAGAT tpg|BK006936.2|:213776-215382 7X257= 303=7X 
 tpg|BK006936.2| 256947 + tpg|BK006936.2| 256898 - INS AAATATTTTAAACAGAACCGGAGATGAAGAACCACTTGTCAATAGACTTGTCAATTGGAGCATCTGCCTTTGGAGAAGCTGGTGGGATGGCATCAGAGGCAGCCTTGGAGTAGGTTGGGGTGTCAGGCAAAGTA tpg|BK006936.2|:256616-257229 7X117= 115S7X 
 tpg|BK006936.2| 119151 + tpg|BK006936.2| 119568 - INS CACTACTTCTTCTTCTTCTTCTTCTGCGTTTATTATGTGCTCTACTGTTGTTATAGTTTTCTATATGTGTGTTATTCGAAATTACCGGAGCCATAGTTTCATTTGTAAGAGCTTCGTCCGCTAATGCGGTGGGTTCTAAGTTCATCATCCCATTTATACCAAATGACGGCCCTAATATAATAG tpg|BK006936.2|:118771-119948 7X4=87S 85S7=7X 
 tpg|BK006936.2| 559932 + tpg|BK006936.2| 560386 - INS GCTTATGTATGTATTATACAAAAGACTTAAGACCTTGAAAGGACCAACCGTTAGGAGCGGATATTGTTAAGAAGTTTATGATGCAACTTTGTAAGGGTATTGCATACTGCCACTCACACCGTATTCTGCATCGTGATTTAAAAC tpg|BK006936.2|:559630-560688 7X5=98S 13S21=1X85=7X 
 tpg|BK006945.2| 900870 + tpg|BK006945.2| 901075 - INS GGGTATGAAGTGTATAGCGTAACAAACCCATGGCTAAAATTCTGCTAACAGGAATGTAATCCTTTTCCAAGCATTTTGCCAATGATGAAACTGTGGAAGATGGGCTACCAGCTTGCTTAAACTTGAAGGTAGCATTAGAGATATCTTGCAGTTCATTGAATATCCATTTTTGAGGTAGTGAGTTTTTCAACATTTCAATATACTGGAAGATCAAGAC tpg|BK006945.2|:900422-901523 7X5=255S 6S198=7X 
 tpg|BK006945.2| 664993 + tpg|BK006945.2| 664777 - INS GACACCCTTAAGATGACATATACAGATGGGCGGCGATAAAGTAAGTTTCCAGAGGTAATACCAGGCAATAAACAGCTTCAATTGCTCGTAACACCATTGTATACCTACAAAAACAGTGGAATAGGGATGAGACATAACTGGCTGGAATTTCAACTGTACTTCTTTGCACAACTAGTCTTGGCG tpg|BK006945.2|:664397-665373 18S23=1X56= 65=34S 
 tpg|BK006936.2| 17498 + tpg|BK006936.2| 17185 - INS GGATTCGTATTACATTTCTGAATGACCATAACATTGCTAGTCTTTTTCTTGAGGGCAGAAGCTCCCCGAATAATATTTTCTTCGACGGCTATCTTTTTTTTAATGTTCTGCTCCAATTGTGAAAAACTCATGACTGTAAACTGCTCCCTATATGTGTGATACTATACTTACTTTTCCTCGCTAGAGCTTCTCTCCGCAGCTACTGTTCTAGGTTTTATTCCTATTGATTATCTAATATAGTTTTAAAAATCTATACTGAAAGGGGATCGACGCTGAATACCTCTAACGTAAGTGTGGACGAGTGGTGGCAGAGACTTTTAC tpg|BK006936.2|:16529-18154 7X248=1X11= 161=7X 
 tpg|BK006945.2| 630469 + tpg|BK006945.2| 630809 - INS GTGCTATCATCAAGTTCATACTGTGCCTGCTTGATCGATAAATGGAATCTCTCTCTGTAATAGCCAATTAAACTGTCAAATGCATCCATTCGCATGGATATTAAGATATCGTCTATATTTGAAATTCTTGACAAGTGCCCGTGAAGGCGCTTCTGTCGGGTACTTAAAATTTCTGGAAATAATGCATGGCAACATATATATCGCAGCCTAGACAACCATTCGTTTAAAAAGGCATTGCTTACACGGGGTGATCCACTGCCATCCGAATTATAGCCACTCAACTCTAAAAAATTGTTCCAAAGATTTAAATAGTTGTCCCACTCGATAGGCGCAAACTCCAGGGGAATGATGAAGTTG tpg|BK006945.2|:629741-631537 7X37=1X217= 335=7X 
 tpg|BK006936.2| 385492 + tpg|BK006936.2| 385176 - INS GTTAAAGGTCGTAACTACACTCAAACATTGGATATAATTGAAAATTTGATGAATATGGCTGGGATGTCACATTGCAGACTCGACGGTTCCATACCTGCTAAACAAAGGGACTCTATCGTCACATCTTTCAATCGGAATCCAGCCATATTTGGATTCTTGTTGAGTGCAAAATCGGGAGGTGTAGGATTGAATCTAGTCGGTGCTTCGCGACTTATTTTATTTGATAATGATTGGAATCCTTCAGTAGATTTGCAAGCGATGTCACGAATTCATAGAGATGGTCAAAAAAAGCCGTGCTTCATATATAGACTTGTCACAAC tpg|BK006936.2|:384522-386146 7X4=213S 300=7X 
 tpg|BK006936.2| 764873 + tpg|BK006936.2| 765043 - INS GTTGTCCTACTGTTAAACCAAGGAACTTCAGTGGGGGTATTGACACCATATTTGAACCGCGGACTTGGCCCGTTTAGTGAAGTGGCGACAAGTTCATTATTGGAACTCGCGGTATAGCCCAACCTTCCATGCTTTAAATAACCCCAACTATAAAACTTTGCATCATATGCCCGTAATTGGTATACTT tpg|BK006936.2|:764485-765431 7X6=87S 88S6=7X 
 tpg|BK006945.2| 695846 + tpg|BK006945.2| 695306 - INS AAATATGGTAAGTACTGCCAATAGTTCTTGTTTCAACTCTTTGACCCTAGCTTCTCTAATGGCAACTTGAGTAACAGCACGGAAACCGTCTTCCATTCTGTAACGGAACGCCTCGACCTGCTTTTGATCGAATTTGTAAGGCTGTAATTCTAATCCAAGTTTGCTCTGTTGTTTGATGATTCGTGAAAGAATCCTTTCATCCTTCTTTGCTGTCTGTAGCATTGATGGCTTATGCTTACCAAATTCTTTCAGTGGGACTACGAATGAAATTGCAGTACCGGTCTTTCCGCCACGAGCAGTTCTACCTACTCTATGCACGTAGGACTTAGCCGTCGTAGGT tpg|BK006945.2|:694612-696540 7X4=194S 5S325=7X 
 tpg|BK006936.2| 28449 + tpg|BK006936.2| 28652 - INS CTAACAAACTTGATATCAGAACCACGTAGAAGAAAAAGAGACTAATAGTAAAAATATCAAGAAAGTTGACCAATTTTTGTTATATATGTCCGTAAAAGTTATGACTTGGCACTGGTCTTGGTTTACTCATCAATCAGCTAGGATCAGCGCTGAGTGACTGCTTGCGGCTGGGCGGCTAAGAAATGGGAATATGTACAGT tpg|BK006936.2|:28037-29064 7X55=44S 1=159S 
 tpg|BK006945.2| 895951 + tpg|BK006945.2| 895208 - INS GTAAACTACACCGGAGATGTCGTCGTTAAGAAACAAACTTAGAACTTGTGAAGACGGTATGTTTTTCAATAGTTTATTCAAATCTTGGTGTCCCAACCCCGTGTCCGTGATATCCTTATGTTTTGTAGCAGAAAATTATGAGTTAGCTTACACAGTGTTACAAACTTACGCGAACTACGAGTTGAAGTTAAATGATCTAGTGCAGTTGGATATTTTGATTCAGTTGTTC tpg|BK006945.2|:894736-896423 7X3=319S 215=7X 
 tpg|BK006936.2| 395124 + tpg|BK006936.2| 395213 - INS CTACTGAATCATCCAAGAGCTCTGCTACATCTTCCGCTTCTTCTAGTGGTGATGCCTCCAATGCTCAAGCTAACGTTTCAGCTTCCGCTAGCTCTTCTTCCTCTTCTTCTAAGAAGTCTAAGGGTGCTGCTCCAGAACTTGTTCCAGCCACTTCATTCATGGGTGTCGTTGCTG tpg|BK006936.2|:394762-395575 75S12=7S 80S7=7X 
 tpg|BK006945.2| 23139 + tpg|BK006945.2| 23589 - INS CCTCAACCCCTTCCCAGCAATCTAGACTATGCTGTTTCTTTTGGCATTCCTACATGGGATTCGGCAATAGGCTATGCGGAAAAGGTGCCAGAGGTAATAGGCAAAATGGCTACAGGATATCCGAGGTACTTTCCTCAACCCCCCGTCCAGAGGCTTTGTGCTTACTTTGTTAAGAAATTTGGGCGAGGTTCAGAAAACTGTCGTCCTTTTCCATCCGTTAACCTGGGTTTAAAGTGTTTCGAGTACGTAAAATCTGTCTCAGGACCTGAAAGTAAAGCTCACCTTGAAGTGGAAACAGTTACGATTAAAAACCGTGGGGCAAAAACGTCGAAAGAACCGGCGGAATTGGTGCTAACCATTGCTGCTGTCCTTGCATCGGAGGAAGAGTTCGAGACTGTGAAAG tpg|BK006945.2|:22319-24409 7X230= 202=7X 
 tpg|BK006945.2| 880545 + tpg|BK006945.2| 880871 - INS GGTTAGTGCATGTTTATTTCCTATTTCCTGTACATTCAGAACGAGAACACAATATATCCAGTTCTATCTGGTTACATTTATGGCAATTCTCGTTCTTACAGAAGTGGATAACTCCCCTGGTTATTTGGCAAGCCACGACGCCCGTTGATGTCAAACCTTGGA tpg|BK006945.2|:880207-881209 7X5=76S 67S14=7X 
 tpg|BK006936.2| 533697 + tpg|BK006936.2| 534139 - INS TTCTACGAGGCTTCTACGAGGTATTGTAGGCCCAATGGTACTGTCGTCCTGGTTGGTATGCCAGCTCATGCTTACTGCAATTCCGATGTTTTCAATCAAGTTGTAAAATCAATCTCCATCGTTGGATCTTGTGTTGGAAATAGAGCTGATACAAGGGAGGCTTTAGATTTCTTCGCCAGAGGTTTGATCAAATCTCCGATCCACTTAGCTGGCCTATCGGATG tpg|BK006936.2|:533237-534599 12S71=35S 107S5=7X 
 tpg|BK006936.2| 185621 + tpg|BK006936.2| 185694 - INS TTTACAGTCTTGTTCTTCTTCTTCCATTACTTTTTTCAGCCATAGGCGGTCATCGTCAGTAACCTCCAGAAGTCTCAAACTGGAAGATTCTTGTAGAATTGACACTGTTAATGGTGAACCGACGAGTTCATCAGTAGATATGTATGTACTGATGGAC tpg|BK006936.2|:185293-186022 7X16=62S 7S1=237S 
 tpg|BK006936.2| 641295 + tpg|BK006936.2| 640604 - INS TTTTTGCTCTAAAAGCCAACTCTAATAGTGCGTAATCTGTGAATTTTTTACCGATTAAAGTAATACCATTTGGCAAACCATCGTCTCGGAACCCTGCGGGAACAGCAAGGGCTGCCAAATCTGCCAAGTTGACAAAATTAGTCCATGTGCCTTGTCTTGAATTGACTAGGACTGGTTC tpg|BK006936.2|:640234-641665 7X3=188S 2S165=7X 
 tpg|BK006936.2| 597493 + tpg|BK006936.2| 597890 - INS GGTCTCAACTGTAAGCAAATATTACGATTATTCTCACTTTTACAAATGAAGAGAAATGACTTAATAGTCACCTCTGAAAAGTGTAATAGCGGAGTTTTCTTCAGCAATTTTAATTATCAACTTCAAGTTAAATCGAATTGTATTGCAAATATTTCTTCTACACTCAGTTTTCTACCCCATCATGAAATAACCGTATACACATCCTTTATTCTCTATCCAAACGTTGTCGATAATATTTGGGAATGCACACGATACGCTATTCAACTTTTGAAGTCCGAAGCAGCACAGTTTACGCT tpg|BK006936.2|:596887-598496 7X217= 148=7X 
 tpg|BK006945.2| 175669 + tpg|BK006945.2| 175698 - INS AAGGATATGATTCAGTAGACGAAGTACAAAGTGGCATATACGAAAAAATGCACAAACAAGTGAATGACACCCCGCATCTACGATTTGGAGTTTGCAGAAGAGAGGCCAGTTTAGAGGCTCCCGTAGGGTTTGATGTGTACGGGTATGGTATTAGAGACATTTCGTTAGAATCTATCCACGAAGGAAAATTGAATTGCGTCCTAGAAAATGGTTCGCCATTGAAAGAGGGTGATAAAATCGGATTTCTACTGAGTCTTCCTAGCAT tpg|BK006945.2|:175125-176242 7X272= 133=7X 
 tpg|BK006936.2| 646580 + tpg|BK006936.2| 646495 - INS GTTTATGTCTAATGGGTATATCATCGAAATTGTAACGAGTAGTAAGGTCTTCATCATTTCTAACATTTTGCGGCGATTCGCTTATAAGACTTTTATTTTCAGAGTCGATCATGGGATAGTCTTCTGCATCCAAGGGCTGATACCCATGTTCATGACGGTCCTGCGCATTTACGTTATTAGTGGTAATAGGAAACTCGAAAGAATTCGCAAGTTTTGGTGAAGACAAAATGGGTTGAACAGGAGATTGAATAGGTGAGTTCTCC tpg|BK006936.2|:645955-647120 7X237= 132=7X 
 tpg|BK006936.2| 590265 + tpg|BK006936.2| 590223 - INS TTTAAGATATATGAGAATATTGATAAGGCTAGAAGGATGGTAGTAAGAAAAGTTGTTGTTGGTAATTTTTCAAAAAAGAGTTTCAAGAGCTGGGAAAAGAATTAAGGCAATGGGAAGCGAACCGTTTCAGAAAAAGAATTTGGGTCTGCAAATTAATTCG tpg|BK006936.2|:589889-590599 7X7=73S 76S4=7X 
 tpg|BK006936.2| 38779 + tpg|BK006936.2| 38965 - INS TCGATTGGACACCACCAAAAATAAAAATTTGAAATCCATTAATTTGGCTATTTCTGCTCGTGGCATTGATGCTCTGAAATCAATAGATCCGGATGCTTGTGAACATATTCTGCAAGATATGATTCCCATGAAAGGCAGGATGATTCATGACTTGAAAGGCAGACAGGAATCACAATTGTATGGCTTGCATGGAGAAGCTATTAATTCTATCAATAGATCTGTATTAAAT tpg|BK006936.2|:38307-39437 7X183=17S 2S1=160S 
 tpg|BK006936.2| 744656 + tpg|BK006936.2| 744687 - INS AAGTTATCCTTTGTATACTAATACTTCTGAAGCCCGATAGACAAGTAAACTTCAATCAGGAGACAGGGGAGAACAAATCTGTACTGGAGGTTTGCAAGAGTCATGGGCTGGAACCCGATCTGCTGAAAAGACTTTTGACTTGGTATACAGAAGAATGGCCTAACAAGAGGTTAAACTCGTTGGAAAAGATATGCAATAAAATCCCAATGCTGAGATTTACAGTATCCAAAGAACTACTGTTGGGCTACTATACTAGTG tpg|BK006936.2|:744126-745217 7X68=1X95=29S 12S1=354S 
 tpg|BK006936.2| 114615 + tpg|BK006936.2| 115173 - INS CCATAGTGGTTGTACAGCAACTGTGATATTGGTATCTCAATTGAAAAAGCTACTAATTTGCGCCAATTCCGGTGATAGTAGAACAGTTCTATCTACTGGTGGTAATAGTAAAGCAATGTCATTTGATCATAAGCCCACATTGTTAAGTGAAAAA tpg|BK006936.2|:114293-115495 7X6=71S 70S7=7X 
 tpg|BK006936.2| 342944 + tpg|BK006936.2| 343490 - INS GCCAGAGGTAAGGATGTCTCTAACGTTTTCATTACTTTCATGAGTGTCATCATGTTTTTGTGGCTGATTGCTTACCCAACCTGTTTTGGTATCACAGATGGTGGTAACGTTTTGCAACCAGATTCTGCTACCATTTTCTATGGTATTATTGATTTGTTGATCCTATCTATCT tpg|BK006936.2|:342586-343848 7X86= 209S2=7X 
 tpg|BK006945.2| 545546 + tpg|BK006945.2| 545130 - INS TGGAGATGAGCATCATTATGTGGTGTTGAAAATATAATATTATGTGGTACTGATTCTGGTAATGTGTATTCTTTCGATATTAGAAACAATGAAAACCGTAAACCAGTTTGGACATTGAAGGCACACGATGCTGGTATCTCCACATTATGTTCAAACAAATTCATCCCTGGTATGATGAGTACAGGGGCCATGGGTGAAAAGACTGTCAAATTATGGAAATTCCCCTTGGATGATGCTACGAACACTAAGGGCCCAAGCATGGTTCTGTCTCGTGATTTCGATGTCGGAAATGTATTGACATCGTCATTCGCTCCAGACATCGAGGTAGCGGGTACCATGGTCATTGGTGG tpg|BK006945.2|:544416-546260 7X4=260S 5S324=7X 
 tpg|BK006945.2| 1010346 + tpg|BK006945.2| 1010991 - INS ATTCAGCAGGATCGAACTGGATTTGGAGTCAGTATTTCCCATTATGCATAGCCTAAGGGAGAATTTTTATGGTTTGATTTGTGTGTATTTCTTTCTCTATTAGCTTTTTCTCTGATTTGTTTGCTTATCTACCTGTACGTGTATGTTGTGTACTCAATAAATAG tpg|BK006945.2|:1010004-1011333 8X129=13S 3S1=166S 
 tpg|BK006936.2| 21511 + tpg|BK006936.2| 21766 - INS ACTACCCCGAACCAAATTCTAAAAGATAGTCAGCTGGATTAGAGTTGTCATCTCCAAACATTAATTTTGCATTATCTTCGGCTTCAATCAAATCGCCTGAGAAGAACTCCTTTAATTCTTCATGAATGTTTGTATGTGGATGACTCTCCATAGTGCCAGCA tpg|BK006936.2|:21175-22102 7X28=52S 1=266S 
 tpg|BK006936.2| 184744 + tpg|BK006936.2| 184990 - INS CCCACTATATAGGGATGTATACAGTCTGGAATATGTTAAAAAATTTAAGACCTTCGAATTATGGCTCACGGATAGATTTTATCCTAGTGTCCTTAAAGCTTGAACGATGCATAAAAGCAGCTGACATTCTTCCGGATATATTGGGCTCTGACCATTGTCCTGTGTATTCTGATTTAGATATACTGGACGACAGAATTGAACCTGGTACGAC tpg|BK006936.2|:184308-185426 21S91= 62=51S 
 tpg|BK006945.2| 788304 + tpg|BK006945.2| 789054 - INS TTTACTACCGACATTGCCTCTCCAAGACATCAAGAAGAAGATATAGAACTTGAAGCCGAACCTAAAGATGCTACCGAAAGTGTTGCAGTCGAGCCATCCAATGAAGATGTAAAACCAGAAGAAAAAGGTTCAGAGGCAGAAGACGATATCAACAACGTTTCCAAGGAGGCTGCCTCTGGTGAGAGTACTACCCACCAAAAAACTGAGGCCTCTGCTTCTCTTGAAAGCAGTGCCGTCA tpg|BK006945.2|:787814-789544 7X119= 165S6=7X 
 tpg|BK006945.2| 132310 + tpg|BK006945.2| 132950 - INS AAAAGCCTGCCTTGTTATTTAATTTGATTAGGAAATTGGATCCAACGGGTCAAAAGAGGATTGTCGTTTTTGTGGCTAGAAAAGAAACTGCTCATAGGTTAAGGATTATCATGGGTCTTTTAGGTATGAGTGTGGGTGAATTACACGGTTCTTTAACCCAAGAACAGCGTTTAGATTCCGTTAATAAATTCAAAAATTTGGAAGTTCCTGTACTTATCTGTACGGATTTGGCCTCCAGAGGTCTTGATATCCCCAAGATTGAGGTTGTTATCAACTACGATATGCCCAAGAGTTATGAGATCTACCTGCATAGAGTTGGTCGTACCGCCAGAGCTGGTAGGGAAGGTCGTTCCGTCACCTTCGTCGGTGAATCATCTCAAGATAGAAGTATTGTACGTGCTGCTATAAAG tpg|BK006945.2|:131476-133784 7X144=1X16= 205=7X 
 tpg|BK006936.2| 340410 + tpg|BK006936.2| 339785 - INS GCCCATATACACCTAGTTGATTTCTGCATTGGCAGTGGTCACGAAGAGATCTTTACCAACAAAACAACAACATGAAACTCTTGGTGTCTGCTCCGGCAAAATGAACTCCTTCAGCAATTTTCCGTTAGTTAAATCGAACATTTGAACCTTACTGGTGGACCAGACAG tpg|BK006936.2|:339437-340758 7X4=174S 147=7X 
 tpg|BK006945.2| 1047235 + tpg|BK006945.2| 1047928 - INS TGAATTCGAAATTTCCCTTAAAGGCGCAAAAAGTCCCTATATGCTTGGCGGCGAATCAGCTGGTTTCATAGTTGGTTTTGATGGTAATGTTAACTTAAAATGTAACGAAGATAATGATCCCAAAAAATTTTTATCCTGCAGCGCAGACAAGGTCCATTTCAGCATTCCCAATTATTTTGCAAAGCCGTTACTGGTATGGTCTAGACCTAGTACCAATACAATGTTCATTCCAAACCAGGACGATACGAACATGCAGAGATATGC tpg|BK006945.2|:1046693-1048470 9S149=47S 59S7=7X 
 tpg|BK006936.2| 489878 + tpg|BK006936.2| 489759 - INS AAGGGAATGGTGAACGTCTGGTTTGCCTCGTTGTATGCCAACCACGCATTCTCGTCGAAATTGATCTCACCAGGATGGTAATGGAATAACGGCCATAGAATAGAATTACTGAACCCGTTGTAGTGTAAGTCTGCGATTTCATCGCTCAGGAAGATGGGTACGGCATTAAACTTTTCCAGCAAGTCCTTCCTCACCTGATCCTTCTCATCGTCAGGAATCTCTAGCCCAGGCCATCCGAACCACTTGAAAGTGTACGTCTTCTTCAACCCTTCCAACGCCGTGACCAGCCCTCCGGACGACATTGCGTACTCGTACTGTCCCGTACTGCTGTTTTTAGTGATTGTCACGGGAAGCCTGTTGGAC tpg|BK006936.2|:489019-490618 7X260= 182=7X 
 tpg|BK006945.2| 914359 + tpg|BK006945.2| 913598 - INS TCTAAGAAGGACATTCTTGAGAATTGCTTAGTTAAAATGTCAAATCTGGCATCAACGTCTGGTATACCAATTTCTACTTCTTGGTCAAACCTGCCAGGTCTCCTGAGAGCAGGGTCGACAGAATTAGGCCTGTTTGTAGCAGCAATTACCACCACTTTACCTGCAGCGCCCATGCCATCCATTAGGGTAAGCAATGTAGCCACGACTCTGCTCTCAACTTCACCGGAGTCATCGTTTGCTCTATTTGGTGCTATTGAATCAATT tpg|BK006945.2|:913056-914901 7X6=152S 132=7X 
 tpg|BK006936.2| 404792 + tpg|BK006936.2| 405359 - INS TTTGTGATGATACTTACGAGTGTAAATAAATAAAAGATGTATTTTGCCAACTTCTCCAATGATCTTTTTTCCTTTGTACATCTAACATAATTGAAGACTTACGAGTGTACATTCACTTTTCATTACTTGGATCTGAAATATTAGAAAGTTACCCGTACCATCAAGAATATAATCGCAGCCCTAATAATTATTCACTGGAGTTAGTCCCAACAAGCATTCCTGTAG tpg|BK006936.2|:404328-405823 7X151= 8S203=7X 
 tpg|BK006936.2| 18329 + tpg|BK006936.2| 18916 - INS CCCTATATGTGTGATACTATACTTACTTTTCCTCGCTAGAGCTTCTCTCCGCAGCTACTGTTCTAGGTTTTATTCCTATTGATTATCTAATATAGTTTTAAAAATCTATACTGAAAGGGGATCGACGCTGAATACCTCTAACGTAAGTGTGGACGAGTGGTGGCAGAGACTTTTACAATGGTTAATAATCAGTCTC tpg|BK006936.2|:17923-19322 7X5=93S 92S6=7X 
 tpg|BK006945.2| 927437 + tpg|BK006945.2| 927982 - INS ATATACTATAAGTAACTTAAAAAGCAACCTTCCTCCCAAACCTACAATCCAATCACGCTGATAAGTATTATCTAGAAAGTTGACAACACCAAGCCATATGGTCAAGAAACATTTATTGAGAGTTATTTTGTAAATAAGACTTTTCGTCATCCATATAAAGCAACCTAATTGTTCATCTAATACTAGAGTCGCTCTTTTGAAAGTTAAGTATAACTACCTCATCATTAGTTGCTACTATGTGTATAAT tpg|BK006945.2|:926929-928490 7X125=60S 1=399S 
 tpg|BK006936.2| 338495 + tpg|BK006936.2| 337910 - INS CTGTTATAATTTTATTTCCATAAATTTAAATTCAAGATTAAACTTCTTTGCTCGTGAAAGTCGAAATTTTTCTTCTTTACTGCTGGCAACATGCACATTCTTTTCTTGTTTATTTTCCACTGTTTGGCATTCAAAGACTTGATTTTTTTTAAGCAATACGTACCATTTGCAGCGGCGGGAGGATATCCCATATCGTTTCTATTCATCAAAGTTCTGACCGCCTCAACGAATTTACTACTTTCTTCTTCCTCTGGAGGGTCCTGGAATAAGTTATCCAAAGAGTCGCAATTACTCAAAGTCATTCTCACACAC tpg|BK006936.2|:337272-339133 7X5=163S 293=7X 
 tpg|BK006945.2| 804936 + tpg|BK006945.2| 804436 - INS GGGTGCAGAGGTAAGCCGCAGAAGACGAGGGAATACTAGGAACAGCGGGTGCTGGTGATAATGGTGCATTAGGAATGGGGGGAGCCGCAACAGATGGCACCGCGCCCGGAATTGGCGGTGCGCTCGCCGATGGAGAGGGTTTAGTGCTTGCATTGTTATTGATATGTTTTAACTTCGGTATACCTCCAGCTAAAATATCGCCCAACTGCGGAGCGCCCATCCCAGGGA tpg|BK006945.2|:803966-805406 7X298= 3S211=7X 
 tpg|BK006936.2| 733085 + tpg|BK006936.2| 733711 - INS CAGCAAATGTTTTCCTGTTTGGTTATACTTGTTCAAAAAACTGTAAAGATCACGTTCATTGGAAACAGATCCAGCAAATGATTTCATAGATTTGGTGGAGTCCAATGGGCTTATTGTAACACCTGTATTCAGAACCAAATTTTCCGTCCATATCGTGTACTTCTGCAATTGGATAG tpg|BK006936.2|:732719-734077 7X7=128S 88=7X 
 tpg|BK006936.2| 732718 + tpg|BK006936.2| 732984 - INS GTTGTTGCAGCAGTGATCCTACTAAATAAATATCCGAATCAGAATGTGGCTTTGATGGTAGAATCATGGAAATGTTTGCGGGATCCTTATCAATTTCCTCCTTCAACTTGCTGACATCAAGTACATTTGCCGATTTTCTATAAATTCCTTCTTGATCAAGCCCAAATTTATCAATAACGTATATGCATTGGCGCACTATCGCAG tpg|BK006936.2|:732296-733406 125S7=1X53= 102=7X 
 tpg|BK006936.2| 412164 + tpg|BK006936.2| 412030 - INS ATTACACATCTGAAAAGCTTCCAGTTATCAAACCTCTTCCATTACACTTAGAAATTCCAGTGCCTTCAGATATTGATATATCAAGAGCTCAGAGTCCTAAGCATATCAAGCAAGTTGCCGAGGAGTTGGGAATCCACTCTCACGAATTAGAATTATACGGCCACTATAAGGCAAAAATTTCTCCAAATATTTTTAAAAGATTAGAATCTAGAGAAAACGGTAAGTACGTCCTTGTTGCAGGTATTACTCCGACTCCATTGGGTGAAGGTAAATCCACTACGACTATGGGGTTGGTGCAGGCTTTATCCGCTCATTTAGGGAAACCATCCATCGCGAACGTTAGACAACCATCTCTTGGCC tpg|BK006936.2|:411296-412898 7X7=13S 180=7X 
 tpg|BK006945.2| 897369 + tpg|BK006945.2| 897503 - INS AAGGACAGAATTCTACAACACCTGTACCTCCAAAAAACCCATTTCTTTTCTGTTTTTACTGAATTGTAATTCGCGCTTGTCTATTCGTCATTCTGAAAAATTTCACGCAAAACAACTGATGACAGATCTTGACCATAGCATAGCATGAAGGTGCAGGAACATGAGGCAGGAGCACCCTACGGGGCACCGCGAAAATAGCTGTGTGAAAGTGCTATGCGATACACATATAATTAATGGTTATTAGATGCGCGCATTTAACATTTTCCCTAACTCAAGTAATAGCTGAAATACCACGAACAAAAGTGTAAATTAGGGTATGTACCAAGTTC tpg|BK006945.2|:896697-898175 7X164= 284S3=7X 
 tpg|BK006936.2| 700490 + tpg|BK006936.2| 700764 - INS GTTCAATATCATGTTCCCGTAGCAATTAAACCATAGGATCCCGAAAATTTTGCCTTGGATAATATCGATCAAAGAGGTGCTGTCTTCTGGCGGCGATGACAGCGCTGCAGTAGTGGTTTCCTCTGCTGACGACATCGAATGACCCGGCGACGGCAGCTGATC tpg|BK006936.2|:700152-701102 7X52=29S 4S1=172S 
 tpg|BK006936.2| 558342 + tpg|BK006936.2| 558763 - INS TAAGAACAGTCTTCAAAGCA tpg|BK006936.2|:558288-558817 7X6=4S 10=7X 
 tpg|BK006936.2| 437217 + tpg|BK006936.2| 437740 - INS TATATTGGTTCAGACCCCCCAATTTTGGAATCTTACAAAATAGAGATAGAAATTAGTCGGTTTTTAAACACAAACTTATATTTCCCCCAAAATTACCATTTAGTCTTACAGCAGTTTACCAAAGTATCCGAAAAGATAAAATCAGTTAAAGAGGAATGTGCCTTACTCTTTATCTCTTATTTGTCTCATAGTATAAGAAGTATTGTTTCGAC tpg|BK006936.2|:436779-438178 10S121=35S 47S6=7X 
 tpg|BK006945.2| 547690 + tpg|BK006945.2| 547598 - INS CATATTTTGAGCTTAAGTACCCTCTTATGCCTCTTTCACTCGCCATTACTGACATTCTGTGATCGCCATTCATATATATAGGCCTGATTGTGCACCAATTGCCGCGCTATCACACCTCCATAAGCGATAGCATTCTTCAGAATATCTTGAAGGCTCAAAACCAAGCCATTGACCGCACAAATCAACTAAAGAACCCATGTCAGACAACGAAAGTTTCTCAAATCCATTAGGC tpg|BK006945.2|:547120-548168 7X209= 116=7X 
 tpg|BK006936.2| 272109 + tpg|BK006936.2| 272211 - INS CCACAGCTCTGCTACACTGCTACATCTAGCGTTGCCGCGGAACATTTTCTCAAATTCCATTGCGTATCAACATCGCCATCTTCATCATCATCATCATCATCATCATCTTCGTTGTCATCTGCATCCTCTCCATTTCCTGCCTCTTTCTTTTTCACAATACGGGGTGCAATGGGCTTGATGTCCTCATCTTTATCCTCCAAGAATGCATCATCATCATTAGAAGCTTCCAGGAGAACGATGGATTCTTCGTTATAGACCATTTTCGATAATAATATTGGCACGATATCCTTAACATATGGTTGTAAGATATGTTCAGGAATATTTGGGCTCGTTGCAAAGGCGTGCAAAAACTCGCAGGCTTCAATAGCCACTTTTTCCTCATTTACAGTGGTGATCAAATGCAACATGAATTGTACAATACCATCTAAATGGGAAACCAGCTTATCTGGTCTGAATTCCAATAAGAAACTAAAACTAATGCAAATCTGTGCCCTAACTAGGTC tpg|BK006936.2|:271089-273231 13S152= 5S483=7X 
 tpg|BK006936.2| 746559 + tpg|BK006936.2| 746606 - INS ATAATGCACAGTCTCATAG tpg|BK006936.2|:746507-746658 7X5=4S 6S4=7X 
 tpg|BK006936.2| 110092 + tpg|BK006936.2| 110099 - INS GGTTCTGTTCAGTATATGAAGTAGCGACAGAAAAAAAGCTTTTATTTCGAGTTCGCATCATTGTCACTTTCCTGCTTTTTCTTGGCGTACTGTCTATCTAAGATAGTCTTTAATATAGCGTCCTCGCCATATTCTTCTTCCTCAATTTTCTTCCATCTCTTTTCTACATCAGCTCTCTTTATTCTACTTTCAATGACAGCACGTTTCTTGTTATTCAAACTTGCCTCCTTGAGACACTTGTTCAAAGC tpg|BK006936.2|:109582-110609 7X8=148S 233=7X 
 tpg|BK006945.2| 105886 + tpg|BK006945.2| 105614 - INS ATAAGTATTATGTAAATATCTAAGCGATCACATGACTGCAAGACCCTTTTCATTGACTTTTCGGTGGTTATGGTATCTCCGCGTTTATTTTTTTCAGGCCATTGTAAGCTTAAAGTTTTTCTGTCGAAATGCTTTATCACCGTTGAATTTAGGTCTGATGGAGAGTTGCCCAATTTATGTTTAGATTTGTAAAACATCTTATCAATAATGTCTGTGGGGAAAGGGGTTCCATTGATTCGTTGCATCATAGCCATATGTTCTAG tpg|BK006945.2|:105074-106426 7X289=4S 247=7X 
 tpg|BK006936.2| 769350 + tpg|BK006936.2| 768891 - INS ATTGGCAATATGCAGAGAATTTGATCTTCTTTTTTGTTTTCCTTCTTTTTTTTCTTTTCTTTGTTTACATAGCACCTGGAACACCCAAGACTTGATTCAAAGCACTTTGACCGCCACTTTGTTGGTATTCAATGGTAATGACTTCTAGCAAAGAAAACCCACCAGCAATGCCAACAACTATACCAGCAGCTTTACCTTTCAAACCCAAAGATTCACCGATAACGGTGATCAAACTTAAGACG tpg|BK006936.2|:768393-769848 7X3=155S 227=7X 
 tpg|BK006936.2| 461355 + tpg|BK006936.2| 460587 - INS TCCCGTACTAAAAAGTCCACTATAAAAAAATGAATCACAGCGTACAAAAGGAAATAACGATAACTGTGATGCTATGTAAAACTATCGTCTTTCCTTTGTTGATAAATATATCCTCAAGGACTACTTCTTTTATATTTCTTGTAGGTGATGTTGTGCCCTCATCGTTAATTTGAATCCCAGCAATTATCAGACAGTTCTGCCGCCCTTCGGCAATGTCCAAGCTGTAGCCAAATACTTAAATCAAGGAACACTAACCATGTATGACATACAAGGAGCACTACCACTGATTTCAACAGATATTAATGGTAGTTTTTTGCAGAATCGTAAGGTAGATC tpg|BK006936.2|:459903-462039 12S40= 168=7X 
 tpg|BK006936.2| 233221 + tpg|BK006936.2| 233761 - INS GTTCTAGGG tpg|BK006936.2|:233189-233793 7X4= 5=7X 
 tpg|BK006936.2| 718107 + tpg|BK006936.2| 718588 - INS TTGTTATTTCTTTTGTTTTCGATTTTGTTATTGTGTCACAAAATAACTAATGGCGACATCGCAGTTTTTTGGGCGGCTGCATACTGTTTAATAAAAAGAAGTTACTGCTACCTCAAGATTTCTTCCTAAGCACTCAAGCCCATGTTTGCCAGTATTGTTATCTTGCAACAAAATCAGACAAATAG tpg|BK006936.2|:717723-718972 7X2=2X25=1X118=16S 2S1=24S 
 tpg|BK006936.2| 147072 + tpg|BK006936.2| 146761 - INS CTCAAGAACTAGGAACGTTACAGTTGGAATTTGCTAGTCAATCGAGTTTCCAATTTCGCAACCTTTATTATAGTACTAATCTTATAAGCCATGGATCGCAAAAAAACACTTATAAACTCAAGTGTTTCTAATAATAACAGTACCATCAAGGGCCTACAG tpg|BK006936.2|:146429-147404 7X233=2S 80=7X 
 tpg|BK006945.2| 41789 + tpg|BK006945.2| 42244 - INS GTAATTGAAGAGTACAATCTTACCAACCACAATGCCCCTTCAGTGAAGGAAATAGCATACGTCAAAGATATACCAGCCATACCCGAATCCAGATTATTAATATTGAATAGAATGAACAAACCAGCTCCAAAAATGACCAAGGATCCAATCATATCTATCCTAAAGGCCAACCAACGATTAGCAACCCACAAGTAGAAGAATGGTTTATTATTTTCATCAATTTTGTGTAAATTCTCTTGCATAAACCTCCCTTCATCACCAAACGCACGAATGGTGGT tpg|BK006945.2|:41219-42814 7X330= 261=7X 
 tpg|BK006936.2| 365645 + tpg|BK006936.2| 366017 - INS GCAAAAGTATCAGGACAGCCCGCACTCTTGCCTTTATCCATTTCTTGCAACCATTCTTCCTGTAATGATTCTGGAAGCATTTGCGATAATAATCGTAAAAGTAGTGTTGAATCTGAATGTGCATCACCCTCACCACTGGTGTTACCAAAGTTTTGAAATAGACCTTGCAGTTGGGATCTGACC tpg|BK006936.2|:365265-366397 7X154=11S 1=202S 
 tpg|BK006945.2| 439114 + tpg|BK006945.2| 439246 - INS CTCGGAAGGAACAACCCATTTAATTCCGTGAAACATCTCGGCTTAAAGTTGAACTCTACCAGTTTCTCGGAAGGAACATGTAAATTTTTGGAGATATACGAGCCCGTTGTCCTAGAACCTTTTGTAGACGTTTTTTCAGTAGAGTTTTTACCACTGTTACTCGGTTGAATAGAATTATGTCGCCTTACTGGAGACCTCAATACGGAAGAATCCGTATCT tpg|BK006945.2|:438662-439698 7X14= 192=7X 
 tpg|BK006936.2| 318634 + tpg|BK006936.2| 318284 - INS GCCCATACATAGTGTTGAGATTGTCTCATATTTTGCATTTTGATTATAACGTTCAGGCCGGTGACTACGTGGCAATCGATTGTACTAATAAACCTCTTTTCGTATTTTTATGGCTTTCTTTGTGGAACATTGGGGC tpg|BK006936.2|:317998-318920 7X154= 68=7X 
 tpg|BK006945.2| 142775 + tpg|BK006945.2| 142954 - INS GAGCAGATGTCCTACATTCATGTTCTTTGTCGAAGGTCTTATAAAGCAGCATGCTCCTGCTGACGAAATTCTTTCATTATTGACAAACAAAAACAGAGGCCTAGAAGAGTTTTTTGTTGAGTTTTTGGTAAGAGAGAACCCGATTAACGGGCATGCTAAGTTTGTTG tpg|BK006945.2|:142427-143302 7X6=77S 80S4=7X 
 tpg|BK006936.2| 568404 + tpg|BK006936.2| 568747 - INS ACACACTTAAACTATCTTTTATTGAAAGACTTGGGATTACAGGATTTACTTTTCCACATATGGCAACCGCTTTTTCATATTCAAGCAACGGAAGACTTACAGTATTCACCGTCAACGGTAAAATTCAACAGGGCGTGGAATAGGATTATATATAAGGACTTTAAATCTTATTTTCCGGAACTGATAGGTACTTTACAAC tpg|BK006936.2|:567992-569159 7X50=49S 6S1=64S 
 tpg|BK006936.2| 346385 + tpg|BK006936.2| 346909 - INS AAATTAGCCCAAGGTTCTATCAACGGTAAAGAAGACTTTTAAAAATACTTTCGTTACATTATTTATTAAAAGAAGAAACGCCATCATTTCATAAAGGTCTCCGGAGGAGCTACTAAAGAAAGAGTGCTGCAATTAATACAATTAATATAAGTGTGGTTATTGAAAATAACTATTCATTTATACGGAGGGTTGGCCGAGTGGTCTAAGGC tpg|BK006936.2|:345953-347341 7X7=97S 101S4=7X 
 tpg|BK006936.2| 480033 + tpg|BK006936.2| 479748 - INS TTAGTTAGCGTTCGTAACCTAGCTTTCGTGGAATACGAGACCGTTGCTGATGCTACGAAAATCAAGAATCAGTTAGGCTCCACTTACAAGCTACAAAACAATGACGTTACCATAGGATTTGCTAAGTAGAATTTCCTTTGCGGAAGTATACCT tpg|BK006936.2|:479428-480353 7X76= 22S4=7X 
 tpg|BK006945.2| 885007 + tpg|BK006945.2| 885724 - INS GTTCTAGGCATATTAAGAAAAAGGATATTCAGACGGTAGTGGACTATTTTTCTGTTCCTGTAAGCAACCCCATGTGTTTCCTGTCACAAGACGCTGCTAGGTCTTTCTTAACTGCTAGTACCTCACAGGATAAGTATAGCCATTTTATGAAGGGTACTTTACTTCAAGAAATTACCGAGAATTTGCTTTACGCCAGTGCTATTCACGATAGTGCACAAGAAAATATGGCTCTGCACCTGGAGAATTTGAAGTCTTTGAAAGCTGAATACGAAGATGCCAAAAAACTGTTAAGGGAATTAAATCAGACTTCAGACTTGAACGAAAGGAAAATGC tpg|BK006945.2|:884327-886404 7X224= 313=7X 
 tpg|BK006936.2| 569597 + tpg|BK006936.2| 570080 - INS GTTCTTGTTCTTTGTTATCTATCATTAAACTAAATAGTTCTGTTGCACTGGTTGCATATTGAAGAATTTGCTGATGTGCACTTGGGTTTGTTATGGCTAATCCTGCGTAAACATGCCACTTGTT tpg|BK006936.2|:569335-570342 7X5=57S 57S5=7X 
 tpg|BK006936.2| 120989 + tpg|BK006936.2| 121109 - INS CTTCTTTGAAACCCGATTAGAGGACCGGATGATGTTATATTTTTGTTAACTAAAGGTGCTATGACTGAAGATTTAGATATTAGTCTTTCAAAATTGAAAAATTTGATAGAATCATACTTAATTCTAACCTTCAACTCCTCGCTGACTTCAATATTAGGTTCAATAATGGGGAAACTTACTGCTCCCATCTTATTGTCC tpg|BK006936.2|:120579-121519 7X118=30S 41S7=1X1=7X 
 tpg|BK006936.2| 64746 + tpg|BK006936.2| 64799 - INS AAATCCA tpg|BK006936.2|:64718-64827 7X3= 1S3=7X 
 tpg|BK006945.2| 590880 + tpg|BK006945.2| 591076 - INS ATTTATCCATTTCTGCATAGATTATTGCCTACCAATGCTTCATTTTCTTTCAAATCAATTAGAAAACAGTGGCAACACAACATGGATATAAATAGTTCGCAAAGTTCATAAAAAGCTCCAATTTGCTCGTCTGCGATACTTGCAAATAGTCTTGTCCTTTTTGAGTACGCAATGAATTGTAAGCACCAGCGAAAAGATTGAAATGCGAGGTTATAATTTTTATCTACATGACCAAATACTCCTTGAAATAATTTTATATATAGTACCAGTTTTAATTTATTCATTGTCTCTGGATCGGCTTTATC tpg|BK006945.2|:590256-591700 24S135= 95=65S 
 tpg|BK006945.2| 421403 + tpg|BK006945.2| 421786 - INS GTATATCTTATAGTCTGTCTGGCATTGTGGAGTTCTTAAGATAACAGAATTTTCTTGTAATTTCAAAAGAGGCCTCATTGAGGTGGTAACAATGTTATCGAATTCGTCAATCTCGAACCAAATCTGCAAAAAAGGGGACGAGGAGGAGCCAGAGGTGGGCGGCACAGGAGTGAAGTTCAGCTGTATGAAGG tpg|BK006945.2|:421007-422182 7X4=204S 96=7X 
 tpg|BK006945.2| 907998 + tpg|BK006945.2| 907678 - INS GACCAGCCTACTGGTGAAACAAAAGTGCTTGAAACAGGTAAGACGTTTATCATTGATATCACCAAAGAAATATATAATGCCGGATTCTATTTTTGAACAGCCCTTTGTTTACTGTGGTGTTTGCCACAGAAGAACATCGCATGGAGATCCATTGAGGCTGACCTCATGTGCTCATATCCTCTGTTCGCAGCATTCTCCATTAACATCAAAGGTGTGTCCTATATGCCGTTCGAGCGATATCTCCATCATTAACCT tpg|BK006945.2|:907154-908522 15S156=1X5= 1S239=7X 
 tpg|BK006945.2| 384468 + tpg|BK006945.2| 384904 - INS CCTTTACATAAAACCGTCACTGTCAACTTTGGAAAAACTAGGATCCCATTCCAAGATGTCAAACCAAGCAGGCATCAATGCACCGCCGTTTGCTGTCACATGAAGCTCTGGAGCATTAGGAAAAACAAAATTAGTATGCTGGAAAGCGGCAGGGTCTCTCTGTTGTAAATACTGAGCTAAAAATCCCCATCCCGAACCTGTATCACCTAATCCATGCAAGAATATGATAGTTTGGCGTGCTGGCTGAATTTTTGCTGCAACTCTAAGTCCATTCATATTCGATAGCGCTCAAATGGGCAAATATAGTGTATGTGTTCTTA tpg|BK006945.2|:383814-385558 7X187=1X24= 160=7X 
 tpg|BK006945.2| 743789 + tpg|BK006945.2| 744534 - INS GTGTGGATTTTAACGAAGTTTATCCGATTGAACCACCAAAAGTTGTATGTTTGAAGAAGATCTTTCATCCAAATATCGATTTAAAGGGGAACGTTTGCCTAAATATTCTTCGAGAAGACTGGTCGCCAGCTCTAGATTTGCAGAGTATTATAACCGGGCTTCTTTTCTTGTTCTTGGAGCCTAATCCCAATGACCCGTTAAACAAGGATGCAGCAAAGTTACTGTGTGAGGGTGAGAAAGAA tpg|BK006945.2|:743291-745032 139S11=149S 121=7X 
 tpg|BK006945.2| 287260 + tpg|BK006945.2| 287641 - INS CCAAATTTGCTAGAAGTGACAGATCAGCAAAAAGAACTTTCACAATGGACTTTGGGTGACAAAGTAAAACTTGAAGAAGGGAGGTTTGTTTTAACTCCTGGAAAGAACACAAAGGGTTCACTTTGGTTGAAACCTGAATATTCAATAAAGGATGCAATGACAATAGAGTGGACGTTTAGAAGTTTCGGGTTCAGAGGCAGCACAAAGGGGGGTCTTGCATTTTGGCTGAAGCAAGGAAATGAGGGAGATAGTACCG tpg|BK006945.2|:286734-288167 7X66=62S 2S1=275S 
 tpg|BK006945.2| 772498 + tpg|BK006945.2| 772391 - INS AAATGAGGAATACTTATTGAACGATCTTATTGCACCTGATGACGAACTGGATATCGAGGAAAACGCCCCTCCAGATATATACTTAGGAAATCTTCCAGAGGATCGTGAGGCTAACGAAAAGGAATTAAAGGAATTGCAAGAATATTATGAGAGCAAGTATAGTGAAGACGCACAATCGGCTGGAACTTCTGGTTTTAATTTAAATGAGGAATACCGCAATGAACCAGTGTATGAGCTGGAATATGACGGACCGGGGAGCTGCATATCACATGTGTCTTATAA tpg|BK006945.2|:771813-773076 7X66=1X256= 265=7X 
 tpg|BK006945.2| 179325 + tpg|BK006945.2| 179751 - INS GCACATATTCTTCGTTCTCCCCTTTTGGAGAGGATTTAAGCTAAGATATATCTTTCTTCGAGCGCAGTGCTGCTTTTGAGTTCTTTCGTTTTAATTTTCCACTTATTTGGCAATAAAAACTGAGTGAAGAGTGCTTCTCTGTCTGTTTTAGGGAGCTTTTTCAGATCATCATCAGATGGGATTTATAGCAAATATAC tpg|BK006945.2|:178917-180159 8X46=51S 1S1=206S 
 tpg|BK006945.2| 725600 + tpg|BK006945.2| 726180 - INS GGGGTCTTGCTGTCGGTGTTCCAGGTGAATTGATGGGTCTCTATCGCCTCTTGAAAGAAAGAGGTAGCGGCCAAGTTGATTGGCGTGATCTAATTGAACCAGTCGCAAAGCTGGGAAGCGTGGGTTGGCAAATAGGCGAAGCACTCGGTGCCACTTTAGAACTTTATGAGGATGTTTTCCTGACATTGAAGGAAGATTGGTCGTTTGTATTGAATTCTACCCATGACGGTGTTTTGAAAGAAGGCGATTGGATCAAGAGGCCGGCACTATCTAACAT tpg|BK006945.2|:725032-726748 7X52=1X32=53S 1S1=172S 
 tpg|BK006945.2| 989845 + tpg|BK006945.2| 989658 - INS CTAAAGCAAGCGCCCTCCCACACGAAAAGAACAATTTGGGGGACATCAATTGCAGTGACGGAAGACGAAAAAGCATCAAAGGAGAACAAAGAATTTCAAGATATGTTATTGCAGCGAATAAGGCAGGAAGATAGTTCGGATGTCACAGATTCGACGGATTCTCCTCCTACAAGTAATGGTAAGCGAGGCAGGAAGAAGAAAGGTAAAGTC tpg|BK006945.2|:989224-990279 7X1=1X83=20S 1=337S 
 tpg|BK006945.2| 737100 + tpg|BK006945.2| 737115 - INS TGTATGGGAGTTTTCCAGAACCGTACAAAATCTTTTCCGCGTAGGTAAATGGCCTGTTTAATCTTTTTCTTACGATATCCAGCGTTTCCACATTCTGCTTGTAGTTAATAAAAGAATGATCTTCTAATAAGTTTTGGTTGACTTTTGAATCTCTAGTCAAGTTGGAGACTGTCGCAAGACCACGAACAATGGGTCTCTTGATGGCAGAACGTGCAGACAGCATTGTATATCTAT tpg|BK006945.2|:736618-737597 7X5=181S 5S215=7X 
 tpg|BK006945.2| 930317 + tpg|BK006945.2| 930550 - INS TTGTTATGCAGTATCTCTGTTAAAGAAAATGATGAATCTTAAAAATTACATTAGTCTGATCGACTGGTTTAATAAAACCTTTGAGTTCAAGCGTTACGGCGAGGATGGATTTGGCATGGGCGTTGAAATTCCTTATAAAGCTAATAGCTGTGTGCAGAGGAGCGCCTCAGTGGTTGAGAGACAAGAATGAATAAATTTTGAATTACAAAAATCTAATAAACTGTGGTACTGAAATTGTATATATTTTCCTATCATTCAAGAGCGTATACTCGTACCCCGAAAGC tpg|BK006945.2|:929735-931132 18S75= 267=7X 
 tpg|BK006945.2| 127310 + tpg|BK006945.2| 127470 - INS GAATGCCAAAAATTATGGTAGTCTGAATAAATTGGCTACTGGTTCTGCAGATGGTGTGATTAAATACTGGAACATGTCTACTAGAGAAGAATTTGTTTCCTTTAAGGCGCATTATGGACTCGTTACTGGTCTTTGTGTGACACAGCCTCGTTTTCATGACAAGAAGCCAGATTTGAAGAGCCAAAATTTTATGTTATCTTGCAGTGATGACAAAACTGTCAAGCTATGGTCAATAAA tpg|BK006945.2|:126822-127958 10S218=1S 9S6=7X 
 tpg|BK006945.2| 1002144 + tpg|BK006945.2| 1002627 - INS AAAATTGATGGGTATCGTCACTTCTCGTGATATTCAGTTCGTTGAAGACAACTCTTTGCTTGTTCAAGATGTTATGACCAAAAACCCTGTCACCGGTGCACAAGGTATTACATTGTCTGAAGGTAATGAAATTTTAAAGAAGATTAAAAAGGGTAAGCTATTGATTGTTGA tpg|BK006945.2|:1001788-1002983 7X6=79S 81S5=7X 
 tpg|BK006945.2| 269917 + tpg|BK006945.2| 270109 - INS ATTCTTATAATTATAATTTCGTAATACGGCAGGAGCACACCTTTTCATAATGGCCAAAAAGCGTGTTTCAGTATACTCCAACACCCTTAATCACTTAAATTCGAAGCTTTGTACACTATTGCGGCCTCTTTCCTGGGTATCGAGGCTGCGTTAGCGTCACCTAGAAAT tpg|BK006945.2|:269567-270459 7X5=79S 80S4=7X 
 tpg|BK006945.2| 672085 + tpg|BK006945.2| 672075 - INS ACCTCCGTCCACGTCCAAGCAACTAAAGAAAAGTGCTTTCCAGATGTCAATGAAGGCAAAGAAATTACTAAGGATGACGCTAAAGTATCTCTCGAGTCCAAAAAAAACAACGAAACTTTTGTTGATTCAAGTGTAGTAGAAAAACATACCCCCCCAGACAAAGACTGTAACAATTGTAACATTACAG tpg|BK006945.2|:671687-672473 7X11=12S 164=3X4S 
 tpg|BK006945.2| 745547 + tpg|BK006945.2| 746075 - INS GGGATACGGTGCAATTGATAATAGGGATAGAGCTATAGTAAAACAGTTTGGCCTAACGGTTGTCTTGTGGGATCTCGATACTTTTGATTGGAAATTAATCACTAATGATGATTTCAGAACAGAGGAAGAAATACTTATGGACATAAATACTTGGAAGGGAAAACGGAAAGGTTTGATCTTAGAGCACGATGGTGCACGAAGAACAGTTGAGGTTGCTATTAAAATCAACGAACTTATTGGTAGTGACCAATTGACAATTGCAGAATGTATTGGTGATACAGACTACATCGAACGCTACGACTAGAAGTAAGATTTCCGAGAAATAAAGTTTCTCTCTATATA tpg|BK006945.2|:744849-746773 7X196= 171=7X 
 tpg|BK006945.2| 797543 + tpg|BK006945.2| 796841 - INS TGTTACAGAATATCATAGCCTTGATCAACAATAAAATCCCAGCAATTATCAAATTATCCATCCATTTCTCAGTGACATTCTCACTAGATGAGCGTTTTTGAGAATAATGCTAACATTTGGTAAGGTATGAAATAAAATGCGATATCCTCCGTAGTTGTCGTCCGATATAGTGTAACGGCTATCACATCACGCTTTCACCGTGGAGACCGGGGTTCGACTCCCCGTATCGGAGATATAT tpg|BK006945.2|:796351-798033 7X4=277S 119=7X 
 tpg|BK006945.2| 550096 + tpg|BK006945.2| 550345 - INS CTCTTCAGTATTGTTATAGTACTCACCCAAACGCATGACCCTATGTAATTTATCCTTTGCAAAAGTAAACGTTTCTTTGTAATTGTGGGATTTATCCTGAGCCATAAATAACTTTGAACCAATGTAGGTGCTCGAAACAGCCAATCTCTTAGCATACCATG tpg|BK006945.2|:549760-550681 7X5=75S 76S5=7X 
 tpg|BK006945.2| 48569 + tpg|BK006945.2| 48723 - INS GTTCTTTTCAGTGTAGTGATTGGCAGTGAAGCTATCCCTCTTTGCCACCCAATTTTGACGGCAGTTCTCATAGCATCTCAAAGCAATAGCAGTGCAAAAGTACATAACCGTAGGAAGGTACGCGGTAGGTATTTGAGTTCGTTGGTGGTTATCCTCCGCAAGGCGCTTCGGCGGTTATTTGTTGATAGTCGAAGAACACCAAAAAAAATGCTGTTATTGCTTTCTCCGTAAACAATAAAACCC tpg|BK006945.2|:48069-49223 16S112= 19=110S 
 tpg|BK006945.2| 1020195 + tpg|BK006945.2| 1020715 - INS GATCATATTGGGAGGAATTTTCGATCATACTATGAATTTTGGTGTTGCCCCTGGGAATTCCAGGTTTTCCATTTCCGTTCATTTCGTTATCTGTTTCTGTAGTGTAATTTTTAGAAAATTCTTGTGTTTCTTGAATGTGGATTTTTCTAATTTTACTGCTCAATTCGCTTCCGTGAGCGCCACGTCTTTTATTTACTGGTATTATTGCTTCATCAGAACTTTCTGAACTAACTTCATCTGTTTCCTCTTCAAGCCCACCATCATCACTCACTTCTGGATTATTTGCATATACAAAATTCTCTCG tpg|BK006945.2|:1019573-1021337 7X245= 5S280=7X 
 tpg|BK006944.2| 534190 + tpg|BK006944.2| 533890 - INS CCATAGATGAACCTTTTCGCTTCTATCATCGTGAAATCTGAGTAGTTTAATTAACAGCGTGTAGACAGCTGTCTTGCTAATGACGTCTTTCCAAACAATCACAGAAGCGACACCTACCAGAGGCCTCAAGAACACCTTAGAACCACATGATGCGTACCTACTACATACAAGGTTCCATCCGTATCTTTCGGTTAACCAGTCGCTGCAATCCAGCCCACTGACTACGCCAATGAACGCTACGCTATCTTCGAAACAAGGACATTCATCAATGGGCCTGACGTGGTTAAACAGAATAAACA tpg|BK006944.2|:533278-534802 7X223= 150=7X 
 tpg|BK006945.2| 129007 + tpg|BK006945.2| 129425 - INS CTCTGGTTCTTTTCTCTGAAGACTACAACCTCGAATAATTTTCCGACTCTTTCCAAAAATTCTTCCACACCAGGTCTTTTAATGACATAGACATTGTGTACTTGGTCATCTATTTCCACAGACAAAACAAAATCCGCAGATCGTAAGTATTTGAAAGAAGAGTGTACCAAGGTTTCATCCAGGTCCAGTATTAGGCATTTCTTGCCCTTTGTACTTTCATCTTGTGGGGGGAGCAGAGTGTTGTAACCTGGTGCATGATACTGGCCCTGCTGCAAAAGCGTTAGATCAATATATTCTTCATC tpg|BK006945.2|:128389-130043 7X29=1X214= 284=7X 
 tpg|BK006944.2| 105181 + tpg|BK006944.2| 104981 - INS ATATAGCTGGAGGTCAATCGAGAAAATCCTATTCCAATTGCAGTACTTGATTCGTACACTCCAAGTACCAACGAACCATACGCTAGAGTTTCTGGTGATTTGAATCCAATTCACGTTTCACGTCATTTTGCCTCTTACGCAAACTTGCCAGGTACTATCACGCACGGTATGTTTTCTTCTGCTTCCGTCCGTGCTTTGATTGAAAACTGGGCTGCTGACAGTGTTTCATCCAGGGTACGTGGCTACACTTGTCAATTTGTTGACATGGTTTTGCC tpg|BK006944.2|:104417-105745 7X4=181S 3S255=7X 
 tpg|BK006945.2| 670703 + tpg|BK006945.2| 671299 - INS GACTAGGAAGAAGAAGAGCAAATCGGAAGGGCAGATGAGCAGAAAGAGGATGAAGAGGAAGAATCTCTCGATGAATTATCCACTCCCATGGTATATCCAATAAAATCATCTATTCCCCATAATCATAACGAAAAGGTTCAGTTAGTCACTCCCGACCGTTCTGTTTCCATAAGAGCTGATGAATGGGATTTAAAGTCAAATACTGAAGACGAAGAAGGTAATGTTCTTGCAGACCTGAAAATAAGCAGCACTAAGGAAACAAAAAGGCAAACAGACTACGTCCATATTGATTCAGAAGACCAGTCACCAGTAGTATCCGCTCAGATGAGAAA tpg|BK006945.2|:670025-671977 13S79= 8=1X157=7X 
 tpg|BK006945.2| 151141 + tpg|BK006945.2| 151491 - INS GTTTAGCCAAGATCCTGTTTTAAGAACTCTAACTTCCTTGGTCCAGTCGCCCTGTATGCTAACAAAAACGTTGTCCAGATGATCTTTTCTGCAGTTTAGTTTTGTACCTAGTTTAGTGCTAATGGAGCCATTGCAGTCTAGTAGGTTTTGCGTTACATTAGCAGGAATCAAATGGAGTTCGAGGAATTTTCTTAAGTTTGTCGAGTTCGCCGTGATGCCACTTAATGGAATAGAAGAAGCCGTTGGAACTAAAAGCGAGTACTCTTCGT tpg|BK006945.2|:150589-152043 18S123= 125=17S 
 tpg|BK006945.2| 274171 + tpg|BK006945.2| 274178 - INS AGTGGACTGGTGGTGGCTTGTTTCTTCGAATGCCTCGACAGCATCCTTAAAGCTATAGCGATGTGTAATGAATGGTTTAAGCGAGAGTTTTCTGCTAGAGACTAGCTCGATGGAGTCACTATAATCACCTTGACAGTATCGGAAACAGCCTTGGAATGTCAGTTCTTTTGTTGGAATGATCGAGATGGGAAATTGTATTTCCTCTTGTCCCATTCCAACTTGAACGATCGTTCCACCTGCCTTACAGACTTCGATGCCTGCTCGAACGCAAGGCTCTGCAC tpg|BK006945.2|:273595-274754 7X4=297S 264=7X 
 tpg|BK006945.2| 1052387 + tpg|BK006945.2| 1052301 - INS GCCCATTATTTATTTTTCCTTTCGTTTTATATGCTTACTTATCCTATTACATTATCAATCTTTGCATTTCAGCTTCCATTAAGTCAGATGACTGTTTCTCAATCTTTATGTCGTCTTTTTATACCGCATATGATAATACACTTGTAACATGAACACTGGTCAATAGATGATGATAGGGTTTCGTTCCAACACCATCACGTTATCAATTCTTTCGTGTCAACTCCTCATTTACGTTATACTC tpg|BK006945.2|:1051805-1052883 7X254= 226=7X 
 tpg|BK006945.2| 761943 + tpg|BK006945.2| 761493 - INS TATGATATATCATCACGTGAGGTGGATTTGATCTTCACAATCTGAGCAATATTGCAGAACGCAAAAATCACTTCCGAAATAGATGATTGAGCTACAATTCGTGGTATTAGGTCCCCATATGTGAGAAAATATCTTGTTGAAGTGATAGCATGAGATAAAGCACTCTTTAAGTATACTATTTCGTTTTCTAAAGAACTTTGCAGTGAAACTGATGATAGGACAGGTAAGAGATCGCCTATCAACTTTGCTATCTTAATTATAGTCTCAAGCAGAATCGGCAGGCGTGTGGTGGTGGTATCCACAGGATCAATTCGATGGAGCGTGTTTTGAAAATAAAGTGTAAATTGAGTTTTTAATGCTCGGAAGACTTCAATGGATATAATACCATTCACGCTCATAAAATCATCGTTTATTTTGAAGGATTCAAATAATGTGTCATTTAAATAGAAATTTAGATCACCCTCGTCTAACCCATTGTTATGCGTCCCCATATCC tpg|BK006945.2|:760489-762947 7X280= 110=1X137=7X 
 tpg|BK006945.2| 230951 + tpg|BK006945.2| 230960 - INS GTATGACCCCTCATACATGCTTGTTCAAACACAAAAGATTGAGGTTGAAAACTTGGCAAGAATTGGGCTAGGAGAAAGTGGCCAGGTGCTTCTTGTTCAGAACCAAGCAGATATGCTAGCACAATGTGCACCGTTCTATTTTTTTCTATAGTGTGTTTACATTTCTTGGCACATTGCGTTCGGTTTCAAAT tpg|BK006945.2|:230555-231356 7X7=16S 96=7X 
 tpg|BK006945.2| 131702 + tpg|BK006945.2| 132397 - INS TAAGAAGAGGAGGAAGCTAAAAAGCAAATGTACGAAAATTTCAACAGTTTGTCTTTATCTCGTCCGGTTCTTAAGGGCCTTGCAAGTTTGGGTTACGTCAAGCCTTCCCCTATTCAAAGCGCCACAATCCCCATTGCCTTATTGGGTAAAGACATCATTGCCGGTGCTGTGACTGGTTCCGGTAAGAC tpg|BK006945.2|:131312-132787 7X11=165S 165=7X 
 tpg|BK006945.2| 781271 + tpg|BK006945.2| 781648 - INS GTTCATTAAGAGCACGTTGCTTGGTCTAGGCCAAGATTACTTAGAAGATCAATATCAAGAGTTCGCAGAACAGCATTTCCAGCCAACCAGGGATCCGTTTTATGAAACGAATAAAGATGGTAAAAAGCACCGCCGCAGACTGCCATATTATTGCAC tpg|BK006945.2|:780945-781974 7X5=73S 72S6=7X 
 tpg|BK006945.2| 79979 + tpg|BK006945.2| 80192 - INS AAGAATCTTTTCATCCATATTACGGGAGCTTTTTTTTTCCACTTAATGTATTGATCTTCCTCCCGTTCTTTGACGATTCGGCGTTGCCCTTAAAACATATGCTTCTATTCCTTTTTTGATCTTACCCATTTATTTGTTTTTTTTTATTTTCCGGTGGACAACAAAATGTTAAAGGAAAAAAGAAAGTACCTTGCTCGTCATCGCGCTTGCATAATGTGCGCCATTACCCTGTAACAAAAACAAAAGATAGAGTGGCAACAACTTGACACAACTTTGCAATTGTACCATGAACCCCAACAAGAAAGGCGGTTGAGAGTAAATGATGTGGTTTGGTTCCTTTTTTTTCCTACATTTAAGGTTCATAGAGA tpg|BK006945.2|:79229-80942 7X365= 184=7X 
 tpg|BK006944.2| 341902 + tpg|BK006944.2| 341905 - INS GCGCTAGGCCACTGTTTATATTTCGCAGTTGTATGGGCCATTTGTTTTGGTGCTATCAATGATAGATCTAAGAGTGCTTGTTTCGAATGGTTGCTAGCATTTTGGTTTGGTATCATATTTATGATTCTTTCCGCCGACTTTTATTTAGGTGGAAGATACAGACAATCCCGCTATTTCAACCACGTGGAATCATTTTCGGGTTATTACAAGTATGACAAGGCGCTAGGCCTCTACCACAGTGAAGACGTTTTGCCTTCGGACGATAACGCCGGCGTGATTGCCACAGAAACAGCATCTTCAAATATTTACAATAATTCCTCTTCCAACGAATCTATTCAAGTAGTCGTATGACCTCATATATGCTAGACTTGACTAGGAAATACCCTCTAACCTGCAAGATATATTCATCTTTTTCTTTCCAAAGCACAATTTAATAAAACTTGCAAGAACATCGTCATCATTTCCCCCTTTTATTTTTGTTATCCCCGTTACTGATGTAACTAATACCTAATTCTATGCTTCTCAATCTGTATAGT tpg|BK006944.2|:340816-342991 7X6=200S 6S514=7X 
 tpg|BK006945.2| 319834 + tpg|BK006945.2| 319351 - INS CTCTGTAGGTTTAGTATGGTAAAGATAATGAACGTCTATGATTTTGAGCAACAATCCAGGAAGAGCTATGTCTCTGTAGGACGGGTCTAACTTTCCTGAAAGCTTTTAACTTTGTACTACTGGCTGAGGTAGAAAAAGGAGTAGTGATATGTGGCATTTTTTCTGCGCTTGAAGTGAGAGTCCTTATATGATATGACTTAATAACGTGAGTTATAGAATTACTCACTGTGAAGTGATTTTTGGCAGACAGTGATAACAT tpg|BK006945.2|:318819-320366 7X144=1X159= 6S237=7X 
 tpg|BK006944.2| 526992 + tpg|BK006944.2| 527279 - INS CCTCTTTCCAAGCTTTTCTTAACGTCCTCTTTTGGTTTTATATGCCCCTTTCCAAGCTGGGTGGATACCCCGTCCATTGAGTGCCCGTGCCCAATCAAGCTAAAGCCAGACTAAAAAGAGGAAGAGTTCAAGAACCATCAATGCCTCCAGCACAATTTCACAACAGCTTGACACTTTGGCAACGGTTATATCAGAGCATAGCGACGGGATTAGAGAGATGCAAGACGACGGAAGAAAGAAGGGAGTGCCCGGCATGCGCTGAAAGCGCCCTGTAGTACAAGCGTACCGCCGTTGAATAGGCCATGGTACATCACACGATGATTGATAATTTGATGCAAGCTGCCATGCTCAGATGGTTGTTTCCCGTTTCTCTCTTTCACTTTTGATCTCCTGCGAAGAATAGGATGAGATGTGAATTTTCGTTTCTAATCCCCTCGGCCG tpg|BK006944.2|:526096-528175 7X304= 414=7X 
 tpg|BK006945.2| 572099 + tpg|BK006945.2| 572005 - INS CTATAAAAGTGGCCATTTCTAGGTCATTGAGAGCCATATCTGTGTCATTAACATGGTAATAGGCCAGGCCACGACGGTACAAAGCTTTGGCCTTGGCTTTTTCGTCAGCCGCTTCGGCAT tpg|BK006945.2|:571751-572353 7X4=180S 60=7X 
 tpg|BK006945.2| 47504 + tpg|BK006945.2| 47509 - INS CCAGTGCTTCTTGACTTCATCGTATTTGTCAGCGAAGTTAGCGTCAATGGTGGAAACCAACTTAGCCAAAGCAGCTTCGTCTTCGGCTCTGACTTCGGTCAAAGCGGCAACAGCAGAAGTCTTTTGGTTAACCAAAGTACCCAATCGAGCCT tpg|BK006945.2|:47186-47827 7X3=73S 72S4=7X 
 tpg|BK006945.2| 604864 + tpg|BK006945.2| 604387 - INS GGTCTCAATTTTTTGCGACAAAGGAAACCTATTGCAAAAAGTGAAGAATGACAGAGAAGGATAATCAGTATATCTCGGTACACC tpg|BK006945.2|:604205-605046 7X55=1X127= 42=7X 
 tpg|BK006945.2| 533018 + tpg|BK006945.2| 532889 - INS GTTCATGGCAAAACCATTCGCCGCATCTTTATATATTTCCTCCACATCCTCAACTTGAGAATCTTCAAGAGGTTTAGCTCTACGAAACCAACTATTGCTTCTTTCTCTAAATCTGAATCGACTCTTTTTCCCATTTTCCGAAGAAGGCACAGCCGAAGTTGGAACATTCAAATATTTTGAATCCTCGCCGTTATTCTTTTGCTCAACTGTAGCT tpg|BK006945.2|:532447-533460 7X365= 1S200=7X 
 tpg|BK006949.2| 310482 + tpg|BK006949.2| 311198 - INS TATATTATACCAAGACTCTGTGCTGTCAACAATTCCTGCCTCGTTTGAACGGTATTATAATCGACTGTCAGGTATTGGGACCTCAAGGGAACTACTACTCTTTAATCCTACAAATGACTGAAAACAATTCAAATTCTGACTACCAATTTTTACTTTTGAATGCTTCTGATTTGACCTCCAAATTGTCGATTAACGGGCCATTACCGGTGTTCAATAGCACCATAAAACACATTCAGCAACCAATCTCGGCCATGAATACCAAGAACTCCAACTC tpg|BK006949.2|:309920-311760 7X293= 8S249=7X 
 tpg|BK006945.2| 643127 + tpg|BK006945.2| 642488 - INS CTCTCTCTTTTATATCTTGTAAATCGCTGCGTTATGTATGCATATTGTACTCCTACCTTCGTAACTGGAAAGAATCAGTCTGAAAGTTTATTGAGCCTGAAACGGAGCAAGATTATAGTTGAATGTTTCTTATTCGGTGTTGATAGTAGATGATGACCAAAGCTTTTTTTAACAAACTACCGTTTGAGGTATTCCGTCGGTACGTTAGGACAGGTAAAAGCATCCCTCAAAGAAGCCCCAGGACAAGAAAATCTCTTCTGGTGGGTGGGACTATTG tpg|BK006945.2|:641922-643693 7X3=319S 259=7X 
 tpg|BK006945.2| 397971 + tpg|BK006945.2| 398119 - INS TCGTTGATGGTTAGGGCTTGGAGAAATTTTTGAAGAGACGTTCTTGCATTCAGGACATGGTATGTTTTTAATTTCGTTTCTTTAGTTCTCAGGCTCTTCAAAGTACTAACACTTTATTGGCAAGGGGCGCTCAAATGTGATGCATCATTATAGAGTAATAATAAAATAAAAAGAAAGGATGCAAGCCCGGAACAAGAGGCAATTG tpg|BK006945.2|:397547-398543 28S49=32S 98S5=7X 
 tpg|BK006945.2| 860758 + tpg|BK006945.2| 860791 - INS GTGAAGGTGGTATTCTATCCGGTGAAATAAAGAATGTCTTACTTTTGGATGTGACACCATTGACATTAGGGATTGAAACATTTGGAGGAGCGTTCTCACCCTTGATACCTAGAAATACGACAGTTCCAGTAAAAAAAACAGAGATATTTAGTACTGGTGTTGATGGGCAAGCGGGTGTTGATATCAAAGTTTTTCAGGGTGAAAGAGGGTTAGTGCGTAACAACAAGTTGATTGGTGATTTGAAACTTACAGGAATCACCCCTTTGCCT tpg|BK006945.2|:860206-861343 7X7=5S 135=7X 
 tpg|BK006945.2| 645266 + tpg|BK006945.2| 645232 - INS TCTTTGCTGACTCTTAACTTTTGCAGCGCCTCTTTGGTGTCGAGTAACTCGTGTTCCAGTAGAACGTTGCGTTCCAGTCGTCGGTCACTCTCCAATTGTAATGTCTCTATCTTATTCCTCAGTTGGATATTTTCATTTTCCAACTCATCTACCTGTATCTCTA tpg|BK006945.2|:644892-645606 7X5=76S 78S4=7X 
 tpg|BK006945.2| 1023888 + tpg|BK006945.2| 1024593 - INS ACACTATTCAGTCTAGAATTAATACAGAATTAGAGGCCTTCGGGTTTTCTTACCATCTTGGAGTTACATGGTTTGCGCTTCTGTGGTGTTTTGCAGGTTTGATTTCTGTGTCATGCTTAGCTTGGTCTGGCTTAGAATGGTGTATTTCCGATAATGGCACGT tpg|BK006945.2|:1023550-1024931 7X1=1X8=71S 40S41=7X 
 tpg|BK006945.2| 428917 + tpg|BK006945.2| 429071 - INS GTTCAAGGCCGTTCATATTGGGCTCCATGTAATATCGGACCATATTCCCAAAGTACTTGGTTAAACGATGATGCAAACCAAGTCAGT tpg|BK006945.2|:428729-429259 7X6=37S 40S4=7X 
 tpg|BK006949.2| 324334 + tpg|BK006949.2| 324630 - INS GCTTACCACCATAGACAGGTCACTTAAAAACGTGGGAACTTCTTGATTCGCTTCATTTAAAATTTCCATCAAACCCTTCACAATATTCTGATTATTACTATTGAAGAATGAAGTAGCCACGCCTGTGTTACCAGCACGGCCTGTTCTACCAATTCTGTGAACGTAGTCATCGATGTCGGAGGGCAAATCATAATTAATGACATGTGTGACATTCGGTATATCCAAACCTCTCGCTGCTACAGCTGTTGCGACCAGGATATCAGCTACGTTAGCTTTGAAAGCAGATAAGGCACGTTCACGTTCAGCCTGTGTGCGGTCACCATGTATGGCTGTAGCTTTGAAATTTTGCATGATCAAAAAATCTGTGAGTTGATCCGCCATTCTTTTCGTTTCAACAAAAATCAATGT tpg|BK006949.2|:323504-325460 7X233= 383=7X 
 tpg|BK006944.2| 179496 + tpg|BK006944.2| 179212 - INS CCAACAGTGGTGAAAAAGGATGTTCTAGTGGTGAAAAAGAGAAGAAAAGAATTCAAAGTTTTCCTCCCATAAGTATACCTATACTTTTTATCTGTGATTGAAAGCTGTATACCAACAGCCTTCTATATATTACCTTGTATACCATTCAGTAGTCTTAAGCATCATCTAACTTTTGACCAGGTCCATTCTGATTGGCTGCGGTAGCCCGCTCCGTTTTCCGCTCTAAGCGTTTGGTACTTGTATAAATGTGCACTGGCATTATGATATCGAGATCCCCGCATAGAAATCTCAGGACCAACCAAAAATTGCCAATCACAAGCTCTAAGAATAATAAACGATGTCTGCAATGATGGTCAAGTTAGGACTGAATAAGTC tpg|BK006944.2|:178448-180260 7X405= 3S361=7X 
 tpg|BK006945.2| 323342 + tpg|BK006945.2| 322859 - INS GGAAACCACTACAATCACAAAAAATACCCCTCCCCTGGCGTGCAAATTCCTGTCAGGAACGCTCTTGGCGAAGTTTCTCCGGCCAAACAAATTGCCCAACTTTTCGCAAGACAGCTGTCTCATATTTACAAGAGCCTCTTCATAGAAAACCCCCCGCTCTCTCCTGAGAACGAGCTGGCATTGACTGCCGTCTTCTATGACGAGACTGTAGAGCGACGCCTTAGAAGGCTCTATATGCGAGCTTGTGCAAGGGCATATACGACTACTAATGCCGACTCCACCACGG tpg|BK006945.2|:322273-323928 7X4=255S 269=7X 
 tpg|BK006945.2| 736455 + tpg|BK006945.2| 736228 - INS ACGTTCAATTTAGCAAAGTCAGCGATCTTACCACGACCAGTTGCTTCCAAATATTCAATCATAGATTTGTTGAATGGGAAAACAGATGTGGTAGCACCGATTTCAGCACCCATATTACAAATGGTACCCATACCAGTAGCGGAGAAGGTGTCAACACCATCACCGAAATATTCAACAATTTTACCAGTACCACCTTTGACAGTTGTGATACCAGCCAATTTCAAAATAATATCCTTTGGAGAAGTCCAACCGTTCATCTTACC tpg|BK006945.2|:735688-736995 7X275= 132=7X 
 tpg|BK006944.2| 68893 + tpg|BK006944.2| 69512 - INS GGTAGAGACGTGCTGGAGCCGGCCGGAGGTAGGATCTTGGTTGAGGCGGAAGATAAAGATCTCTTGCTGTTGGTTGTGTGAGCGAAAGAGTTTGCACGGCGAGAGGTTTTCAACGAATTCGGCAGTTTTGGGCTGGAGGATTCGCTGTCATTAGTACTTGTAGAGTGGAAGTCTGGAGGTAGAGACGCCTTTTTCTTCAACTTGTTCCCAT tpg|BK006944.2|:68457-69948 13S33=66S 68S14=31S 
 tpg|BK006949.2| 899619 + tpg|BK006949.2| 899827 - INS GTGTGGACCGTCACAAACGAGAGGCGGCGGGCTAGTCGTCGCAAGCGACAAATCTCAACTGACAGTAAATAACGGTGATAAAACAAAATTAGCGCAATCTCTCAAACTACTGAGGACAACCAACTTGAATTGCACTCTTCCAAGTTGTAGCATGGCTTGGGGGGTGTGTGATCCCATCCTGTATTATGGCAAAGCAGGCAAAACAACCGCTCTGCCGTCCGGGTAACTTTTCTTGTTCCACCTCTTTTCCCCAACATATATGAACATGAGATGGTAAGAGCAAGAAACAACGGTTCTATGAGCAACGCAAAAACAGCACAGCACACACAGCAC tpg|BK006949.2|:898939-900507 7X158= 313=7X 
 tpg|BK006944.2| 597699 + tpg|BK006944.2| 597913 - INS TTGTACCAATATCATGCTACAGTCTACACAAAGTATAGCCATATCTGCTTGTGATATCCCCATTATAGCGTTTGGAACAAAATCTCTATGGCCTGGCGCATCCACAATAGTAAAATTTGCCCTATGGGTAGAGAAATGCGATGTACAAATTGACACTGTTACACCACGTTCGCGCTCTTCATTTGTCTGATCCATAATCCATGCAAATTTGAAGGATGACTTACCCATAGTTTCACTCTCTCTTTGTAGCTTTCTCAGTTGGGATTGGTTGACAATGTTCAGATCATAAAGT tpg|BK006944.2|:597101-598511 7X5=180S 274=7X 
 tpg|BK006945.2| 937662 + tpg|BK006945.2| 937940 - INS TCATTTTTGGAGATAAGGTGATTCTAGATGAAAGAATAGAGAATTGGCCAACTTGCGACTTTTTGATATCTTTCTTTTCTTCAGGATTTCCCCTAGATAAAGCAATTAAATACGTCAAGTTACGCAAGCCTTTCATTATCAATGATTTAATAATGCAAAAGATTTTGTGGGACAGGAGATTATGTCTACAAGTATTAGAAGCCTACAAC tpg|BK006945.2|:937230-938372 7X174=15S 1=41S 
 tpg|BK006949.2| 883754 + tpg|BK006949.2| 883814 - INS CCTGCGTAACCCTATTGCACATACTGATGACAGGGAAAAATGTGGAAGGTTGCGACAATTTGGCCTACCGACCTGCGTACAATTATGAAATGACGTTTTCTCCAAAGAAGACTCATTACTCATTAAGTGAGCTGAATCTCGAACGAATAACGCCAAGGCCGGATTTGGAGGGAAGTGCCTCTCAAAAAGAAAAAAAATTTTTAATTTCTGAAGAAGATTATTTATTATTGCAGAAATTGAAAGCCTCTCAAACATATAATGATTCCAATGCTGACAAAAATTTGCCTTCCTTTGAAAAAGGTCCTCGTATGCCCAGTCGGGGTCGACCCAGACCGAGAGAGAAGGAAATAATCACCATCCAATATGATTTTGAATTACCAGGAAGAGCCGATATAC tpg|BK006949.2|:882948-884620 7X202= 12S47=1X324=7X 
 tpg|BK006945.2| 293355 + tpg|BK006945.2| 292601 - INS TGGCTATAGATTTCTCCTTATAAACTCTGTTAAAAAACTCAGCTATCATTTGATGACATAATATAGGTCTCCTTTTACTTGCTCTCTTTGTTGTGTGGAGCAAGAGGGCCCAATATATGACTGTTAACTTTTCACAAAGACTTTTTTCTTTATTATTGGAC tpg|BK006945.2|:292265-293691 7X4=160S 141=7X 
 tpg|BK006945.2| 998875 + tpg|BK006945.2| 999646 - INS TATAAGCAAATGGTCGTAACAACAGGGTGGCTTCTCATAACCAAAATTTCAGCGCTAGTATATACGACGATCCACAAGTTTCGCAAGCAAAGCAGACGCAGGTACCGGCTGCTATTACAAAACACAGAAGTTCAAATAGTGTTTTATCCGGTGGTTCTTCGAGGATCCTGACTGCTTCCGATTACGGTGAACCCAATCAAAATGGACAGAATGGAGCAAATAGGAC tpg|BK006945.2|:998409-1000112 7X7=5S 113=7X 
 tpg|BK006945.2| 141720 + tpg|BK006945.2| 141105 - INS CTATACTCCGAAAGAATCTCCGAATGTAAGAATGATGCTTCGTAGGTCTATGTACAAACTTTACAGCGCAGCTGATGCAGAAGAACATCCAACTATCAAGTATGAAGACATTAACGATGAAGATGGCGATTTTACCGAGCAAAACAATGATGTATCATAC tpg|BK006945.2|:140771-142054 7X69=1X129= 80=7X 
 tpg|BK006945.2| 226368 + tpg|BK006945.2| 226801 - INS CATACAAAATCAGAAATTTTATATTCAGCCGCCTTTTTCTCATTTTTATCCTTGCTGTTGTCATTATTGTTATCACCATTATAATCATCTTCGTCAAAATATGTAGCGAATAGCAGATTCCCAAATTCTGTGTAAAAATGAATGTTAACACTATCC tpg|BK006945.2|:226042-227127 7X4=74S 73S5=7X 
 tpg|BK006944.2| 284004 + tpg|BK006944.2| 284294 - INS ATATTTTGCATAAACTTGATTCTTCTCTTCTTATTTCATGTTTCAGTGGGGCATTTTCCATTGTACTTTTGCAACAATAGCGAAAAAAACAATTTTCCGTAAAGAGAAGCGTCAGTCATAAACGGTGTATGTTACCCGAACTGGAATGAATTTTATCTTAAGACTGGAAAACAATTTAGGATAGAACTGAAGATAGTGCAACACGTCTGGTGATATCATGTGCTTTCAAGCAGGATTTGTCACAGTGCTTTAGAA tpg|BK006944.2|:283480-284818 7X135=56S 1S1=163S 
 tpg|BK006945.2| 1060846 + tpg|BK006945.2| 1060779 - INS CCTATCCCAGAATATGGTTAGAAAGATCTTAAGCTAGATAAAGAAAAAGAAAAAAATAGAAAAAAGCCTGCCCGCTTTATAAGAACTTTTCTCAATATCTGTTGAGGAACACTTAGTAATATCGTCTATCATGGTTGCTTTATTCTTAGTGATATTACTCTCTGGGATTC tpg|BK006945.2|:1060425-1061200 26S194=1X21= 149=7X 
 tpg|BK006945.2| 795611 + tpg|BK006945.2| 795912 - INS GTGTTGAGTTACAATGATCTTAGCGACCTGTGCTCATTATTTGCTCCACTAATTCTAATTTTCCTCGCCTTTCATATTTCGTATCTTTATTCTATATCCTAAAATTTTTTTGGCAAATCCCAGATTTGGCTTTGATTTTGGCATCGGTTCGGTTCTTTCAAATATCTTCTTCCCGTGAATCAACTGCAC tpg|BK006945.2|:795219-796304 11S158=9S 14S4=7X 
 tpg|BK006939.2| 116970 + tpg|BK006939.2| 116486 - INS GTACAATTTTTTACTCTTCGAAGACAGAAAATTTGCTGACATTGGTAATACAGTCAAATTGCAGTACTCTGCGGGGGGTGTATACAGAATAGCAGAATGGGCAGACATTACGAATGCACACGGTGTGGTGGGCCCAGGTATTGTTAGCGGTTTGAAGCAGGCGGCGGAAGAAGTAACAAAGGAACCTAGAGGCCTTTTGATGTTAGCAGAATTGTCATGCAAGGGCTCCCTAGCTACTGGAGAATATACTAAGGGTACTGTTGACATTGCGAAGAGCGACAAAGATTTTGTTATCGGCTTTATTGCTCAAAGAGACATGGGTGGAAGAGATGAAGGTTACGATTGGTTGATTATGACACCCGGTGTGGGTTTAGATGACAAGGGAGACGCATTGGGTCAACAGTATAGAACCGTGGATGATGTGGTCTCTACAGGATCTGACATTATTATTGTTGGAAGAGGACTATTTGCAAAGGGAAGGGATGCTAAGGTAGAGGGTGAACGTTACAGAAAAGCAGGCTGGGAAGCATATTTGAGAAGATGCGGCCAGCAAAACTAACTCGAGTAAGCTTGGTACCGCGGCTAGCTAAGATCCGCTCTAACCGAAAAGGAAGGAGTTAGACAACCTGAAGTCTAGGTCCCTATTTATTTTTTTATAGTTATGTTAGTATTAAGAACGTTATTTATATTTCAAATTTTTCTTTTTTTTCTGTACAGACGCGTGTACGCATGTAACATTATACTGAAAACCTTGCTTGAGAAGGTTTTGGGACGCTCGAAGTCTTCCGCTTCCTCGCTCACTGACTCGCTGCGCTCGGTCGTTCGGCTGCGGCGAGCGGTATCAGCTCACTCAAAGGCGGTAATACGGTTATCCACAGAATCAGGGGATAACGCAGGAAAGAACATGTGAGCAAAAGGCCAGCAAAAGGCCAGGAACCGTAAAAAGGCCGCGTTGCTGGCGTTTTTCCATAGGCTCCGCCCCCCTGACGAGCATCACAAAAATCGACGCTCAAGTCAGAGGTGGCGAAACCCGACAGGACTATAAAGATACCAGGCGTTTCCCCCTGGAAGCTCCCTCGTGCGCTCTCCTGTTCCGACCCTGCCGCTTACCGGATACCTGTCCGCCTTTCTCCCTTCGGGAAGCGTGGCGCTTTCTCATAGCTCACGCTGTAGGTATC tpg|BK006939.2|:114116-119340 7X72=3I484=30S 849S9=1X7=148S 
 tpg|BK006945.2| 432662 + tpg|BK006945.2| 432171 - INS TCTATGAGATGGATAATGTGATACGATCTATGGAGCAAGAATATCGGTTAATATTGCTCTTGAACCATAGGAACAAAAATCAACATAGAGCGGCTAGCTGGTATGGATCGTTCAATGAGATGAAAAGAAATTGTGGACAAATAATAACGCTTTTTAGCTCGAGAAGATTACAAGCCAAACGCCTTAAAGATGTTGAATGGGTCAAGTTGCACAGGCTATTACAGAGAGCACTTTTTAGACAGTTAAAGAGATGGTACTGGCAGTTCAATGGCGTAATTGCGCTGGGACAATTTGTAACGTTGGGTTGTACACTAGTAACATTGCTGGCAAATGTGAGGGCACTGTATATG tpg|BK006945.2|:431457-433376 7X5=276S 175=7X 
 tpg|BK006945.2| 618473 + tpg|BK006945.2| 617805 - INS GTTGAAGCCCACTGATAACAAAGATCAAGAAAATTTGAATAAATATTTTCAGGGTGAATTCACGAGACTCCCTTGGCTTGACGAAATCACTATAAGCAAATTAAGGAAACAACGGGAAAATAGGACTTGGCCTCAGGGCACCTTTGTCTTAAACTTAGAATTTCCAATGTTAGAGCTTCCTGTTGTGTTCATC tpg|BK006945.2|:617405-618873 266S12=28S 181=7X 
 tpg|BK006945.2| 678879 + tpg|BK006945.2| 679153 - INS TGAAGAACAACTCTTTAAGATCGCTCACTGTCAAAATCATACGTATTGAAAAATGTTCATCCATCCGAATCCAGGGATTTTACCTACCAAATCTGCAGGAACTGTTCATCAACAATACCCTTTGCGACACCACCCAACACCAAAAACAAGCGTCAAATGATATGAGTTGTATAGAGTTCACTT tpg|BK006945.2|:678499-679533 7X4=87S 88S4=7X 
 tpg|BK006945.2| 679972 + tpg|BK006945.2| 679947 - INS ACGTGTTGTACTACAGAGAAGATGGGCTGCCTCTTTGTACGTCTGTGGACAACGAAAATGATCCCTCATTATTTGAACAAAAGCAAAAGGTGAAAATCGTCGTTTCCAGATTGACACCACAGTCTGCCACGGAGGCTACTTTGGAAAGTGGCTCCTTTGAGATCCATTATTTGAAGAAATCCATGGTGTACTAC tpg|BK006945.2|:679545-680374 17S87= 68=36S 
 tpg|BK006944.2| 142935 + tpg|BK006944.2| 143656 - INS GATTTACGTGCCACCGAGTAGGTTTCTAAAATGTGCAACCATTTTAGGTATGTGCGCAGCTCTTTATTCTAAACGGGAGTCACTACATTACTATTATCGTGTTTTTGCCCATGTACTTTCTCATAATCTTAAGACAACAACGGGATGATAGGCGCATTCGGACTTTCATTGATGCAAATGTGTGAAAAATGCATCCAAAAGACAACTTTTGTACAGAATACAATTGCAAAAATACTTTACGGGCATAGATCGGTAAGGTCACCGGGAAGCTAGCGTAAGAGACCTTATTCGGAACCGAGCAACCATTTCCGAATGTAGTAGTAGTTGAAGGAGTAAATCGACCTTATTGTACACTACTTCCTTTAAATTTGATTTCTGGCCC tpg|BK006944.2|:142157-144434 7X328= 191=7X 
 tpg|BK006945.2| 437356 + tpg|BK006945.2| 437530 - INS TTTGAGGTGCGGAATTTGACGACGAAGTTGCGATAGAATCAGCAGCAGGTGTGCCAAGACTTGCGTTAACATTGTTATTAGAATAATCGGCGGTTGGTGCCGAAGTCGATACTCTCCTTACCCTGAATGAACATCGTCTCTTGTATGGATGAGCTACGTC tpg|BK006945.2|:437022-437864 7X5=75S 77S3=7X 
 tpg|BK006945.2| 157974 + tpg|BK006945.2| 158586 - INS GCTATCATGAAGGAATAGTTCTTTAACTTGCTGCTTCTTAAACTTCTTTGTTTCCAGGCCAGTTTGGTTAGCTCTGATATGCTCAACAACTTGAATTTTTTCCTCTTTGTTTAGGAACCAAGCATTGGTGACGTTATCTGGAAGGTATAAGAATGTTAGAACACCAAACGCAACTGTAACCAGACCAACGACCAAAAACATTATTTGCCAAGAGGTGAAAGCGGTACCATGATAATGTAAAAAGCCAAAAGAAATTAACCCGCCCACAATATAACC tpg|BK006945.2|:157408-159152 7X9=149S 138=7X 
 tpg|BK006945.2| 816629 + tpg|BK006945.2| 816619 - INS CCCGTGTTTTTTTCGGAATTCGGCTGCAATCTTGTAAGACCAAGGCCATTCACTGAAGTTAGTGCCCTTTATGGCAATAAAATGTCCTCTGTTTGGTCTGGTGGCCTTGCATACATGTATTTTGAAGAAGAAAATGAATACGGAGTTGTTAAGATAAATGATAATGATGGAGTGG tpg|BK006945.2|:816255-816993 7X93=38S 1=198S 
 tpg|BK006945.2| 122118 + tpg|BK006945.2| 122339 - INS TTGTTCTAGGGCTTGTTGCAGGATTTTTGCAAATCGAGTCAGTCCATGGGTTTATTTGGTTCCTGATTCTGTACAACTTGATTAATGTCATTTACATTGTTTGGATCTGTCAACTTAAACCAGGAAAGTTCTACCAAAGCCCACTTCATGACATTTTTTTCGAATCGTTTTTTAGAGAGATAACTGGTTTTGTCATGGCATGGACATTTGGATACGCCCTAATCGGAT tpg|BK006945.2|:121648-122809 7X5=109S 111S3=7X 
 tpg|BK006945.2| 136892 + tpg|BK006945.2| 137366 - INS GCGTATGATAGCAAGCTTTTGATTGTGCACTCGTAAGTGACTTGACTGGCTTTCCTAATTTAGGATTCAGTAGCAATTTTATGTTTTCCAAGCTTTCATCTGGCATCTGCCTGTTATGCTTCATTGCTTATGCCGTTATTTGAGGTTACTTTAATCTATTTTCCTACTGATGACACAATTGAGTCAATCCAACGTGGAACGGGTTGCCCTTGTATACATTTCAGTTTA tpg|BK006945.2|:136422-137836 7X4=110S 108S6=7X 
 tpg|BK006944.2| 108327 + tpg|BK006944.2| 108718 - INS CGCGTGTCTATCATCCAAACACATTACAACATCCGTACATTTAGTTGGCTCCATTTTTTGAAAAAATACTTCCGAGTAAGATGCTGAAAGTAATCAAATTCCGTGAAAAAGGAACCGATTTGGTAAGGGCGGACCTGCCGGAAGAAAATCGCTCCCGCGTGTCTAC tpg|BK006944.2|:107981-109064 7X10=10S 146=6X1S 
 tpg|BK006944.2| 327517 + tpg|BK006944.2| 327925 - INS TGTGATAGTAGCCCGAAAGAGTTATACCGAAAGGTAACGGTACTGGTGGCACTGGCGTACCGCCGTTATTTACAGAAGTTGGAAGGCTGGTATTGTTGTTCAAGCCAGCGGTGCCAGTTGGATCCATCAACTTCATTTTCTTAGTTTCTGGCTGGTTGCCATCTTTAGAGCTTCCGTGTAGTTCCTCTTGTTTCTTCAAAAACGTTTCGACCTCCTTTTCCTTGTCCTGGTCGGGTACTAAAGAATCGAGAAGGATATCGCGGGTTTCGCAATTGGGGCATACAA tpg|BK006944.2|:326933-328509 145S14=1X76= 5S263=7X 
 tpg|BK006949.2| 902333 + tpg|BK006949.2| 902461 - INS CTGTACTTGAAGTCCATCGCTTTACAAAGTGTTGTATCGAAATGGCTGGGCTCTGACTGGGAGCCCATCCTATCGAAAATTGCCGCGAAAAACTACAATATGGTACATTTCACCCCTCTACAGGAAAGAGGCGAGTCTAACTCGCCTTACTCTATATACGACCAATTGCAGTTCGACCAGGAACACTTTAAGTCTCCTGAAGACGTGAAAAATTTAGTTGAGCATATACATCGCGATTTAAACATGCTTTCATTAACAGATATTGTTTTTAACCACACAGCTAATAATTCTCCTTGGTTAGTTGAGCACCCGGAGGCTGGGTATAACCACATCACTGCGCCACATCTAATCAGCGCCATAGAGCTCGACCAAGAATTGCTCAATTTTAGTAGGAATTTGAAATCCTGGGGCTATCCTACCGAACTGAAAAATATAGAAGATCTCTTCAAGATCATGGACGGTATTAAAGTGCATGTTTTAGGGTCGTTGAAAC tpg|BK006949.2|:901333-903461 7X481= 247=7X 
 tpg|BK006945.2| 1004135 + tpg|BK006945.2| 1004135 - INS TGGTATGTTAGCGTTTCATTCAAACCTTCAGTCCCACGAGCTAGAGCACCACGAGGTAAGACACCGGCATTCATAGTTTTCAAATATTCCACTTTTTCGCTCTCTTCTCTTAGCACCGAAAACATTCTTGAAACTTTAGCAATAGCTAATATCTTATTTCTCAAAGCCTTTCTTCGGGTTTCATCTTCTAATATCGCTGATGACGCCTTTTCATCAGAT tpg|BK006945.2|:1003683-1004587 14S107=50S 51S4=7X 
 tpg|BK006945.2| 516561 + tpg|BK006945.2| 516478 - INS TTGTATACGATTTATGCTCTGCTGCAGCAGGTTCTGATGGTGCAGAAGGGCGCGTAAGATCCACTTCTTTCTTCACAACTTGTTGTTCGTCTTTTGTTATTGCATCTTCGTTCTTGTCGACGGTCTGTTCTTCTTCGTTTACGCTATCGGCATCATCAATAAATTCAGGTACCTC tpg|BK006945.2|:516114-516925 7X96=35S 1=173S 
 tpg|BK006944.2| 132892 + tpg|BK006944.2| 132152 - INS GCATGAACTTCTTGCAAATAATTTTGTAAACTTTTATGAATTCTGCTTGATAATGAATTAATCAACTTCAACTCATCACTGCCCAATGATGCGTCGGGATTCACTATTTTTAGATAATCTTCCCTTCCTTGCGTGGGCGAGCTGCGGTTGCTATCGTTAGGACTTTGACCGGTTCTTTTCTCATGGTTTGTCTGAGATTTTTCTACGTTTGGCAGAAGAGATAAAGCGTTTTCAATATCGCATTCATTTTTATGATGTTTGAATAGACCAGAAAGAGTAATACCTAATCTTGGTCTAGATAATGATCCCTGTCGATGTGCCGGTAAGGAGTTACCTTTCTCTAATTTCGCAATTACCCCTGATAACTTTATATTATGTTCATGACTTCCGTCTTCGTAAACTTTGAAGCCATTTTGCTCAATTATACATTGCACATCTGCTCCTGCAAAT tpg|BK006944.2|:131238-133806 7X5=91S 436=7X 
 tpg|BK006945.2| 137855 + tpg|BK006945.2| 137846 - INS ATCCTTCATTCCTTGAATGATTTTATTGGAAGAAAATCACCCGATCTGCCTGAATATTTGGATACCATAAAAATAACTGAACTGGATACAGGTGATGATTTCCCCATTTTCTCGAATTGCAGAATACAATATTCGCCAAATTCAGGAAATAAAAAGCTAGAGGCTAAAATTGATATAGATTTAAATGACCACTTAA tpg|BK006945.2|:137440-138261 7X4=94S 92S6=7X 
 tpg|BK006949.2| 129998 + tpg|BK006949.2| 129906 - INS GGATCAGGACTCAATGTTTGCCCACTAAGAAACCACATTACAAGCCATTACTGCTTTCGCAAAACGCACTTGATGAGTTTAATTTGGTGCAGGATCAGGACTTGGAGAAAATACTATCCGGTGAGAAAGTATATTATTCCGATAGTATCTTTCCCTATAGTACAGTGTACTCCGGATTTCAATTCGGCTCATTTGCTGCACAGCTGGGAGACGGACGTGTGGTAAACTTGTTTGATCTTAAGGACAAGTGTAGCGGACAATGGCAAACGTTTCAGTTGAAAGGTGCCGGTATGACGCCATTTTCTCGGTTTGCAGATGGGAAAGCT tpg|BK006949.2|:129240-130664 21S149= 153=17S 
 tpg|BK006944.2| 9572 + tpg|BK006944.2| 9959 - INS CTTCCATGGCCCAATGCCAGTACACCACTTCTGTCTGCCACATATCGAGCAACTTGAACTCTACGAGACTTGAATATTATATTTTCAGGATCGTATTCATAACCGTATGCCAAAAAAACGGTATGAAGCACGAGATATCCAAGAATAATGATACCCTCTAATCTTGTAGGT tpg|BK006944.2|:9216-10315 7X7=78S 81S5=7X 
 tpg|BK006944.2| 418084 + tpg|BK006944.2| 418167 - INS GAATAACGAACTATAACTCTAAACTGCTTAATGTCAGGAGAAGGACTAAAGAAGAAGCAGAGAAGGAATTTATTACCATGCTGAAGGAAAATCAAGTAGACTCTACTTGGTCATTCAGTAGAATTATTTCAGAACTGGGGACCAGAGATCCAAGGTATTGGATGGTCGATGATGACCCCTTATGGAAGAAAGAAATGTTTGAGAAATATCTTTCCAA tpg|BK006944.2|:417636-418615 7X11=97S 103S6=7X 
 tpg|BK006945.2| 753681 + tpg|BK006945.2| 753938 - INS GCATATGTGTATGGGTCAATATCCAAGAGCTTCAATTTCTTCAATCTAAAAAACGCTGAAGAAGCAGAAGATGGTAAAGAAGACGAAGACATGTGTATCGGTGATTTATTGTCACGTTTAGTTGTCTGTACGACTGCCGATACCGAATCTTGTTGCTTAGGAT tpg|BK006945.2|:753341-754278 7X5=76S 77S5=7X 
 tpg|BK006945.2| 335883 + tpg|BK006945.2| 336305 - INS CTTTAAAAGAGATAACGAACTTTCTGCATTGGAACCGTATCTTACATAATTTACTACACTGATGTAAACACCTTCGAATTTAATATATGGCCTTTCCCTTAACATACGATAATCATCACCCCGCCATATTTCCTTTTCAAAGGTATTTATATCGGTGATTCCG tpg|BK006945.2|:335543-336645 7X37=44S 7S1=8S 
 tpg|BK006945.2| 294665 + tpg|BK006945.2| 294984 - INS CTGGTATCATTTCCTTCGTCTAGCATCAATGGGCTGCCAGTCGTTTCACATGTACCTGGACTGGAACGTTTTATGGAAACCGGTTCGACGATAACACCAACTACACGATAGTTACCTTCACCACGATCGTGATATTCAATCATAATATCGAAATGGTTGGCAAAGTAAGGCAATTCGTAAGTTTTCACCATGTTACGATCATTACGTGTTTCCAATTCCACATCC tpg|BK006945.2|:294201-295448 11S165=27S 24S5=7X 
 tpg|BK006945.2| 436663 + tpg|BK006945.2| 437136 - INS TAATACGGTATACTACAGATCAAAAAGTTCATTGTTTTCCCCTGTGGCCACTGTTTTCACTGGAACTGTATAATCAGGGTAATACTGAACTCAAATGATTATAACTTGAGGCAGAAGACGGAAAACTTCTTAAAGGCCAAAAGTAAGCATAATTTGAATGATTTAGAAAATATCATTGTAGAGAAATGTGGATTGTGCAGTGATATCAACATCAATAAAATTGATCAGCCAATATCTATTGATGAAACAGAATTAGCCAAATGGAATGAATAGTAGTATTCTTTTTTAGTCAGGCTGAAAC tpg|BK006945.2|:436047-437752 7X5=156S 283=7X 
 tpg|BK006945.2| 568988 + tpg|BK006945.2| 569371 - INS CATTATTATTAACAGGGCTTTCTATCTATTCGGAATAAGAAATAATCCCTTCATCCCTATAACAGGGCTTTCCTTTTCTACATTTAATTTCTATCATAAATGGTCTGCCTACGTTTGTTTCATGTTGGCCGTTGTACACTCAATTGTCATGACCGCCTCGGGAGTGAAAAGAGGTGTGTTTCAAAGTCTGGTTAGGAAATTTTACTTTAGGTGGGGTATAGTGGCAACGATATTAATG tpg|BK006945.2|:568498-569861 7X12=76S 6S218=7X 
 tpg|BK006945.2| 311105 + tpg|BK006945.2| 311486 - INS CTGGTGTTCTGTCTTTGAATTACTTCTGGTGTTCTGAATAGAATTAAAAGAAGTGCAAACCTCTTGAATAAGATTTCCCTGGTCACTACAGTACTCAAACAGCCATTCCATTTGAGATTCGTCTATGGTAATATCTGATGACGTTAAGTTTAATGAGTTAACTTGTCTATCTTCTGTAGAAGACCATACTTCGAAACCCTCAATCCCTAGCGACAGTGCAGGGGGACGATCTTCAGACAAGTCTGGATTTTTCTTCTGGTTAACAGTCACTCTGACAGTTTTTACCTTTGCTAAAGCTGCTACTTCTAATAATTTATTTGTTCGGTTCTTCTCTAGAGACTTTTCACTCATTTGATAATCAATACGATCTAAATAGAGCTCAAAACCTTCCTC tpg|BK006945.2|:310305-312286 7X217= 197=7X 
 tpg|BK006945.2| 820735 + tpg|BK006945.2| 821061 - INS CATTTGGACAAGGACAGAAAAGCTTTGATCCAAAGAAAGGGCGGTAAGTTGGAATAAATTATGTAATTCCCTGAAAACTTCCTCGAAATTTATTGCACTTTTTTTACTCAAACCATTTAATAATCATATGTAAAACGTATAAAATAGTATCCATTCCAC tpg|BK006945.2|:820403-821393 7X5=74S 75S5=7X 
 tpg|BK006944.2| 145684 + tpg|BK006944.2| 146454 - INS TAAGCGATTAAGCCCATTTGCTTTTTGTCGCACCGTTTAGGTTCGCGTTAGCAAGATGGAAAAAAAAGAACGCGAATCATGTATTGACGTATGACGTATTAGGCAATTTACAAGATTAAACTTAAATTTGCGACGGAGTTTTGAAGTAGAACGAACACCTTACTCA tpg|BK006944.2|:145338-146800 7X8=75S 76S7=7X 
 tpg|BK006945.2| 261407 + tpg|BK006945.2| 261672 - INS TTTCTAGAAAGCCTGGAGTTGATCAAATGTTCAAAAAATAGGGCAGAATAGCATAACACACATCAATAACACCGAGCCAGCATGCCTACCGTCTACGTGAACAAGCAGCAATTATTTGATCTTCTAGGCAAAAACTACACTTCCCAAGAGTTCGATGAATTATGTTTTGAATTCGGTATGGAAATGGACGAAGACACCACA tpg|BK006945.2|:260991-262088 7X4=46S 45S106=7X 
 tpg|BK006945.2| 26438 + tpg|BK006945.2| 26247 - INS CTGTAAATCAACTACTCTCGAGACCTAATTTCGGGGTGATCTTCTTCACCTTTAGTTGACCAACGTTTTCTTTTGCAAAAAGGTTTGAAAAGTTACCGTCAGCTCTCAAAGCAGGATCATGGTATTCGTGAAATTCCAGCGGGCCATACTTTTCAGTAGGATCCCATGTAGGCAAATAATCTGGATACTTCGATTTCTCTCTATAAGATTTACGGATTTTCAATAAACCAGATGGAGAGACCTCATC tpg|BK006945.2|:25739-26946 15S112=1X79= 232=7X 
 tpg|BK006945.2| 411777 + tpg|BK006945.2| 411237 - INS CGGCGCTCTATTGACTTGAACGTCCCAGCCAAGTTATTGGAAACTCCAATTGACTTGTCTTTGAAGCCAAACGACGCTGAAGCTGAAGCTGAAGTTGTTAGAACTGTTGTTGAATTGATCAAGGATGCTAAGAACCCAGTTATCTTGGCTGATGCTTGTGCTTCTAGACAT tpg|BK006945.2|:410881-412133 7X4=148S 150=7X 
 tpg|BK006945.2| 373129 + tpg|BK006945.2| 373125 - INS ACTGTGGCAGAAACTTCTCCTTAAGAAATTAGGAACTCATAAAAGGAATCAGCAGCTCTATGTAATATCAAAATCTTTTCTATTTTTTGTATTTATGCTCTCATTCATTAATTCTAACGGAGCTATTTATTATAAACAGTGAAGATATAAACCATATGTCTAATAGAACAAATTTCAAAAAGTCTTCAATTTCGTGGATGTGGGAATGCATTTATTAAAAATAATGAATGGCAACATACGACACCAAAATAGGAACACTTTCAGTACTATACAGAAC tpg|BK006945.2|:372557-373697 7X230=20S 6S1=283S 
 tpg|BK006945.2| 793091 + tpg|BK006945.2| 793396 - INS AAACATATAAATGCCTGAACAATTAATTTGGATCCGAGGTTCCGCGCTTCCACCATTTAGTATGAATCATATTTATGTAGTATATAGGATAAGTAACATTTCGTAAATCAAGCTGATAATCCATTTTGACAACTGGTCACTTCCTCAAGACTGCTTATATTAGGATTGTCAAACCACCTTACTATGAATTGCGTTTTGACACAGGAAACGCTAATGTAATATAATCCGTGATAGTTTAATGGTCAGAATGGGCG tpg|BK006945.2|:792569-793918 7X225=13S 2S1=211S 
 tpg|BK006945.2| 121257 + tpg|BK006945.2| 121340 - INS CAATATGTACGGTATTGG tpg|BK006945.2|:121207-121390 7X3=6S 5S4=7X 
 tpg|BK006945.2| 445341 + tpg|BK006945.2| 445097 - INS TGTAAATAGCGGCACCCAGAGAAAGGGACATCTTGGTTCATTTATTGTAGTACTAGAAAATCGTTTCCACCATATAAAAATGATAGACCTTGATCAGACACATGTAGAATTACCGATAGAAGAAATACTATATGAGTACTGTAACTTGTTTTACCTCTTATACGTTACA tpg|BK006945.2|:444745-445693 7X8=34S 46S81=7X 
 tpg|BK006944.2| 482081 + tpg|BK006944.2| 482284 - INS TAGCAAATCATCTTTGTTTCGCGTCGATGCATTGGTATTTTTCTTTGAATGGTAAAGATCTTCATAATGCGAATTATCCTCCTTTATTGCTTGTTCGCCATCAAAGGTAATGTCGCGCTTAGGAACTTTTTTAAACTTTATTGGTTGTAATACACAAATGTCGTTGTCATCATCTTCAGAATCGTTCGACACTAGGGGCT tpg|BK006944.2|:481667-482698 7X6=94S 95S5=7X 
 tpg|BK006944.2| 576397 + tpg|BK006944.2| 576696 - INS CTTCCTCATTGTCGCACAGGCCCAAAGCAATTTTTGATAATGTGTTTGCAGTTAATGGAGCTACTACCAGTATATCCGCCCAGCGACGTAGTTCTATATGAAGTACAGGATCAGTTCGTTGTTTCCATGCGTCCCATTCATCTTGGTCGGTCCATAGTTGAATATGTGGGGGTAACTCGACTACTTGAGCCATGTTGCATTGTCCTGGTGTTGGTGTCACTGGAGTTGCCGGAGTGGATTCGTACTGCGACATTTTATTTAGTTTTTCTGAAGATTTGATAATTTTCTTGGTATATCTTTGTTCGAAAAACTGTGTTGCTGATTGAGTGAGGATAACTTGAATGCTTATTCTATCACGTCCATATATTTCTTCTAGTTTTTTAATCATTGGCTTGATCTTAAATACCGATAACGAACCTGTAGCGCCAAACAACACGTGCAATTTTCCATCATCTTGAGGT tpg|BK006944.2|:575461-577632 7X229=1X79= 231=7X 
 tpg|BK006945.2| 355709 + tpg|BK006945.2| 355889 - INS CAGCCGCAGATAATTCAATATACGTCAGTTCGTCAATTTTACCATGAGTTGATTTTTCATTGATTAATTTGAGAGCGTTCAAAGAGTTGAGTAGCAGACGTAAACTTGATAATAAGTATAACGACTCTGGAGATTTGATCTTATCTGAATACTTGCTGAC tpg|BK006945.2|:355375-356223 7X4=76S 77S3=7X 
 tpg|BK006949.2| 35462 + tpg|BK006949.2| 35487 - INS CCTATATACAAGGATAAAGTGGTGAAAGTCACCGTAGAAAACACACCGATAGCAAAGGTTTTCCAGACTCCGCCAACAAAAATCACGACACCTAATAGTCAAGTTTGGGTCCCTTCGACAAGAAGAAGAACCCGATTGAGGCCTCCCACCCCCTTATCACAGTTACTTTCACCAAGAGAAGGGCGTTTAGATAAAACCC tpg|BK006949.2|:35050-35899 7X4=95S 17S14=76S 
 tpg|BK006945.2| 211595 + tpg|BK006945.2| 212207 - INS GATTAGTTCAGCGTACGCATAGTTTAACGTATATTTTATAGCGCTTAAACTTGGGCGGGCATTAACCTTACCGTATTTCTTCAAATCGTAATCGTGCAATCTTGGTTTAACAATGGATGAGCCCAAGTATAATGAATGAGGCATCACAGTGGCACCTAAGATACCCAATGAAATGTAAAGAGCTTGTTGTTCCAACGGGGAAAAGGAAA tpg|BK006945.2|:211163-212639 11S189=2S 7S7=7X 
 tpg|BK006944.2| 163429 + tpg|BK006944.2| 163620 - INS GAATGAGGAACAATCGTGATATTATTATGTAGAAATATCGATTCCTTTTTGGGGATGCCTATATCCTCGAGGAGACACTTCCAGTATATTCTGTATACATAATATAACAGCCTTTATCAACATTGGAATCCCAACAATTATCTCAAAATTCACCAACCTCTCATGGCGCATATTCATCATGCATGTAACTACCACATCAATGTTCAA tpg|BK006944.2|:163001-164048 7X3=291S 104=7X 
 tpg|BK006945.2| 916330 + tpg|BK006945.2| 916449 - INS ATCATTGGGGTCTATGGTTTGTAATTCCTCTTGTAATACTTTGATTTGTTTTTCATGTTCAGGTTGTAAAGTTTCTTTGGCATTCTCACTAAAAGAATACTTGATCATTTCTTCAACTCTCAACGCCTCAATTCTTAAAAGATTTAATATCATATTGTATGTTAATCTAAACTGAGACTGCAACCTCGTCGGAACACCCATCGTTACTTCTTTGAACGTAGCAATAGATAAAGGACTATTATATGC tpg|BK006945.2|:915824-916955 7X5=46S 231=7X 
 tpg|BK006945.2| 162903 + tpg|BK006945.2| 163350 - INS CTTTTGGTATGGAAACTGTTTAGGACTAGTAGAGTATGGTCTTTGCGGGCTTAGCATTGGCGCCTCGTTGGGAGGAAAATCCACATTGGTAGTCGCGGCCACTGTCGGCACGGCGGCAAAGGCGTCGTATAATGCTCCTCTTTTCTGCGTAGGTTTAGGATGCTGGAGAACATTCCTGTCCTTTGCAAGGTCTTTTGAAAGACCAAATGATCCTGCTGTGGGGCTCACTGAACTCTTGGTATTGCTATTAACGGAAAGGTTGGCGCCACTTCCAGCAC tpg|BK006945.2|:162333-163920 7X8=52S 261=7X 
 tpg|BK006945.2| 1016761 + tpg|BK006945.2| 1016786 - INS CGATTCTTCTTCA tpg|BK006945.2|:1016721-1016826 7X1=5S 3S4=7X 
 tpg|BK006945.2| 580627 + tpg|BK006945.2| 580700 - INS GCCATCAGCACCACAACTGATCAGTTGTTTTTGCTTATTAATAAACGAACATCTTTGAACCGCATTGGTATGACCTTCCAATGTTTTCATAACGCTGAATGTATCCAATGACCATATCTTGACTGTTTTATCACCTGAAGAAGTTGCCAATAATTTATCATATTGGCAAAATGATACATCCCATAGTCCACGCTTGTGGTTG tpg|BK006945.2|:580209-581118 7X6=95S 96S5=7X 
 tpg|BK006944.2| 624811 + tpg|BK006944.2| 624844 - INS GGATTACCTACAAATCTGTTAACAATGTACAAAATCCATTACTAGGATTACCTAGGAAAATCGAAGAGAATTCAAATTCACCATTCAATCCGTTACTTTCCGGTGAAAAACTCTTAAAGCTAAATTCTAAGTCTTCATCAGGTGGATTTAACCCTTTTACCTCGCCATCCCCAAATAAGCACTTACAAAATGATAATGACAAAAGGGAGTCGTTGGCTAACAAGACAGATCCACCAACTCATTTGGAACCCAGCTTCAAC tpg|BK006944.2|:624277-625378 7X158=1X169= 244=7X 
 tpg|BK006944.2| 215198 + tpg|BK006944.2| 215066 - INS CATTATCTCCTCACGTCATAGAGGCCAATTCCTAATGATGAAAAATGAACCTGTAGTTTTCACGGGAAGTGATGATCATTGGTTTTATACCTGGAAAATGCAGTCCTTTAATCTTTCAGCAGAAATGAATTGCACTGCTCCGCATAGAAAGAAACGGCTGAGCGGCAGTATGAGTTTAAAAGGGCTGTTGAGAATTGTATCTAATAAGAGTACGAATGATGAATGTTTGACAGAAACGTCAAACCAAAGCAGCTCACACACATTTACCAAC tpg|BK006944.2|:214510-215754 14S185=45S 29S5=7X 
 tpg|BK006945.2| 414868 + tpg|BK006945.2| 415156 - INS CATTATTGATACCATCAGAGAATGGGCCGATGTTCAAGGAATATGTCTGAGAAACGATAAAAAGTAGTGCCGAATGATTGAGAATTTGACAAAACAAAAACAAAACAAAACAAACGTTACGTATAGATGAAGAATACACGTACACAAATATGCATATATAC tpg|BK006945.2|:414532-415492 17S22=48S 73S8=7X 
 tpg|BK006945.2| 302775 + tpg|BK006945.2| 303224 - INS AGTAGAGACTACTTCGAATAAAGACCTCGAAGATGAGAAGATGAAATTTCAAGAATCTTTGAAAAAAGTGGATGAGATTAAAGCACAACGTAAGGAAATAAAAGATCGAATATCATCTTGTAGCTCGAAAGAAAAGACCCTGGTTTTAGAAAGAAGAGAATTAGAAGGCACCAGGGTGTCTCTAGAAGAGAGAACAAAAAATTTGGTAAGTAAAATGGAAAAAGCAGAAAAGACTTTGAAAT tpg|BK006945.2|:302277-303722 7X8=7S 227=3X4S 
 tpg|BK006945.2| 415299 + tpg|BK006945.2| 415695 - INS TCTATACCGTCGCCA tpg|BK006945.2|:415255-415739 7X3=4S 4S4=7X 
 tpg|BK006945.2| 1048793 + tpg|BK006945.2| 1048841 - INS TTGCCGAATTTGCTGGTTTAAAGGCTAAATCTTCTCATTTTATTATGGATCTTCATCAAAGGAAGGAAGTATTGACTGAATATCAAGCCGGCTTGAACGTCAGAAGGAGAGTTATGAAATTAAAATTTCTGGCTGGTGATGTTGTATGCCAGGACGTGGACATCCGGAC tpg|BK006945.2|:1048441-1049193 7X62=22S 10S1=8S 
 tpg|BK006945.2| 644539 + tpg|BK006945.2| 644121 - INS GTCGAGTAACTCTATGAGAGGCGTATTAATCAATTGTATTTTTATGATTTTGTGTTGTGGTGGAAAAAATTTATTCCGAAGACTTGGTTGTCATCTTAAATCGTTAGCGTTCTTTCTACTTGTAAATATATACGTAAAATTATATATAACAATTTTATATGTGTCATTAAACGGAAGACGTTGTTGCTATCACAGTGGAT tpg|BK006945.2|:643707-644953 7X175= 175=7X 
 tpg|BK006945.2| 154149 + tpg|BK006945.2| 154542 - INS ATAAGATAATTCGATGTCTGCATCAAGACAGATATAAGGTAATAGCGCGTAAAGCCCATCGACGAATTTGGACAAATCCACATTAACTTTCATATATTGTGTATTTGAAATAAGTGAGAATGCACTAACGATACAAAGCAAAGCCTTACGGACCTCAGC tpg|BK006945.2|:153817-154874 7X97=22S 3S1=13S 
 tpg|BK006945.2| 426083 + tpg|BK006945.2| 426324 - INS GCTCAAAGGGATCCCAAGTGCTCGTTACTAATTTGCTAAAATCTACCCAAGACAACTCTTATGCCAAATCGAACATTGTGTTGGGGCAATTACTAGGTATGGCAGATAATGTTACCTATGACCTAATTACCAACCATGGCGCTAAAAACATAATCAAGTATGTCCCATGGGGCCCACCATTGGAAACTAAAGATTATCTTTTGAGAAGATTGCAAGAAAACGGGGATGCTGTGAGATCTGATA tpg|BK006945.2|:425583-426824 7X13=4S 3S225=7X 
 tpg|BK006945.2| 91892 + tpg|BK006945.2| 91286 - INS GACTCCATCTCGTCTTG tpg|BK006945.2|:91238-91940 7X1= 11S5=7X 
 tpg|BK006945.2| 538638 + tpg|BK006945.2| 538164 - INS AAGGAGATAAAAAGACGGAAGAAAATTGAGCATGTTGATGATGAAACGCGTACACACTAGTGCATCAATATTTGCACACATATATTCGCATATATATATAGTAAAATCTAAAGTAATGTAAATATTCCAGGGAGAATCAGCAGAAACGAGACGAAGTACTTCTTAACAAAAAGCCAGATAAC tpg|BK006945.2|:537786-539016 7X5=1X5= 91=7X 
 tpg|BK006945.2| 408192 + tpg|BK006945.2| 408478 - INS CTTATAGAAGTTACTCGGTCGGTTACCAAGCAAGGTCCAGATCGAGTTCTCAAAGAAGACATTCGTTAACACGCCAACGTTCCTCGCAAAGACTGATTAGAACCATCAGTATCGAGTCTGATGTGTCTAATAT tpg|BK006945.2|:407912-408758 7X10=149S 67=7X 
 tpg|BK006944.2| 3520 + tpg|BK006944.2| 4052 - INS CTTTCGTGTCAGGCATAATGACTTAGAAGATAATTTGCTGTTGTCTAATTCAAAATAGGTCTCAAGGACATTAAAGCACAAATGTAATGAATTTAGTGGAGCCAGGACGCTAAAATTGAATATTCTCGCATCAAAATCTTGATGTGTTAAGGTATAAAGATTGGATAAACTTCCTATCATATGGAGAGTTGCATGCCATAATTGAAGTTCGGTGAACTCATTACCATTTAAATTAGATGCATTTAAGTAAAAATCCAACGGCTTAAACATTTTAATGGTGAACTTTTTTAAGTCCTCGATGATGAGTGGAATGTCAGGCGGTTTCTCACGAGCATGAATTTGTTTCATAATATTTCTCAGTCTTAATGTTGTTTTATACAGAAGGATGTCCCCTGATGAAGAATAGTTTTCTAGACGTACCTTGTTTACAAAATCGTCGTTGATTCGGACCGGAATTCCTGTAGAGAGTGAAATTTTAACGTCCGTGAAT tpg|BK006944.2|:2526-5046 7X5=159S 475=7X 
 tpg|BK006949.2| 760162 + tpg|BK006949.2| 760931 - INS AAGGGAAATGGTAATACAGCAGTTAGAATTCCATTTGGAAATGTCATACTGACGTCAGATATTTTACTATTTTTACTTGACAATGTACCTTTACGGAGAACGAAGGTATCTTCCATTTTGAACATTATAAATCCTTCAGTATTCCTCACTATACATCAAGTACTGGAAGTTCTTCATTTAGTGGACAAATTCGATAGCCCTGAGACCTCATCATGTACTAACACAAACGACAGATCATTAAATATTTTAGATTTAGATATTGATCGATTGCCCAGTTTTAACTTTGAACTACTAATGTCGAATTTTATTTCAAGGCTGCATATATCAGATGAGGAGAATGTGACGTTTAAGGTCTTCAGCACACATGCTCTCTTTAGCCGTAACAACTTGTCTATGACTCCTAAAAAGGGACAAGTAATGCAAATACGTCCGGATTGGCCATTTGCGAAGACAGCCCTAGTATCTGATCAATTATCTAACTATATTAAAATTGTGGGTACATCACTCTCTTACCTGAGAATTCCAACAGAGCAGGACGCTAACCCAGTGTCTATACC tpg|BK006949.2|:759034-762059 7X166= 279=7X 
 tpg|BK006944.2| 152974 + tpg|BK006944.2| 153620 - INS ATCGAATATAGATGAAGAGGAGGTAGACTCGGACGAGGAGAGGATAGGCCAAGTTAAAAGAGGCAGAGGCGCCTTGGTAGATAGTGACGATGAATAATCCGGTCCTGAGAAAAAACCATATTTACTTAGGTCATATATATTTTATATTTTAAAGCAACCACCCGTAAGCATTTAAGTCTCTTAAGCCAACAAATCGCCTCGCCATCTTAATCATCGTCATCAGTATCGAATATAGATTTTGGTGGGAAAGCGGTTTTAACGTGGTCCGCTAATTGCATCTGTCCATTTCCATCGTTCGTGGGACATCTATCAATGGTAATTGCGCCCACCTTTGATTTCAATAACGTGAAAGTACCATTGTTATTTTTGTCTGGATTATTAGGCAATAGTTGGCTAGCTTCCAACCGCTGCTGCTGGTCCTGTTGTATATGACTTTGTATATGCCTTTGTGGCGCATCCTCACATTTGCTGAAATCGAATTCGGGAGGTGGTGATGCTGGGGGCGATATCAGGAACATTTTTTC tpg|BK006944.2|:151912-154682 7X4=199S 508=7X 
 tpg|BK006944.2| 622055 + tpg|BK006944.2| 621353 - INS GTACTATCACAGTTAACCGAAACTAAGAGAGACCTCGAATCTCAAGTACAAGACTTGCAAACTCGTATCTCGCAAATTACTAGGGAGTCTACTGAAAATATGTCACTTTTAAACAAGGAGATACAGGACCTGTATGACAGCAAGAGCGACATATCCATTAAGCTTGGAAAGGAAAAATCATCGAGAATATTGGCAGAGGAACGATTTAAACTACTTTCGAATACGTTAGATCTAACTAAAGCTGAGAACGACCAACTG tpg|BK006944.2|:620823-622585 7X4=330S 242=7X 
 tpg|BK006944.2| 123989 + tpg|BK006944.2| 124604 - INS ACGTAAACATTGACGTTATGAAAAGTCAAATTATTCCGCTAATGAAAAAAGCCTGTTACGTTGGCTTACTGACAGCAATCCCAATTTTATTGGAACCCATCTATGAAGTTGACATCACGGTCCACGCCCCCTTGCTGCCAATAGTAGAGGAACTTATGAAGAAGAGACGTGGAAGCAGGATATACAAAACAATAAAAGTGGCAGGGACACCATTGTTGGAGGTTCGTGGACAAGTTCCGGTTATTGAATCTGCAGGATTCGAGACAGATTTGAGATTATCTACGAA tpg|BK006944.2|:123403-125190 7X192=22S 1=284S 
 tpg|BK006949.2| 24475 + tpg|BK006949.2| 24810 - INS TGTTAAGCAACATCAAGAGGTATCAAAGTTGCAAATCCCGTGTGGTCTACTATTCCATTTATTAGCGAATCATTTTGGTCTGATGAGTCATCTGCTAACAGAAAAATTGTCAAAGAAATGTTCAACGATTTCTTGAATGCTGGCGCAGAAATATTGATGACTACAACATACCAAACGAGTTATAAATCAGTTTCTGAAAACACCCCAATCAGAACTTTATCCGAGTACAATAACCTTTTAAACAGGATTGTCGATTTTTCTCGTAATTGTATTGGCGAAGACAAATATTTGATTGGCTGTATTGGCCCATGGGGTGCTCATATTTGTCGTGAGTTTACAGGCGACTATGGTGCTGAGCCAGAA tpg|BK006949.2|:23735-25550 15S358= 341=7X 
 tpg|BK006944.2| 217123 + tpg|BK006944.2| 217360 - INS AAATTAAGTAAACAAGATAAACAAATTGAAAAAACAGCCGCCCAGAAGATATCGAAGTTTGGTTCGTTTGTGGCTGGTGGGCTAGCAGCATGTATAGCTGTTACAGTTACTAATCCGATCGAATTGATTAAAATCAGAATGCAGCTTCAAGGTGAAATGTCAGCATCAGCTGCAAAAGTTTATAAAAATCCAATCCAAGGTATGGCGGTAATTTTCAAAAACGAAGGTATAAAAGGTCTGCAAAAAGGGTTAAAT tpg|BK006944.2|:216599-217884 7X26=1X112= 240=7X 
 tpg|BK006944.2| 161513 + tpg|BK006944.2| 161437 - INS GTGTTTTGGAAAGTGGCGGAAAAAAATAAGAGATATGGAAAACAAATATGAACCATCATTAAACTTGAAAAAGATGAGAAGAAAAGAAATAGTTAGGCTTTAAGTGTCTGTATTGATCAATTAATTATTACTTTACCACTGCTGTTTATTAGCATAATAGCACACGGGATCAGAATGCTTAGTAATACACTTATTATTGCCTGTTTATTGGTGATAGGGACAACCATAGCGCTAATAGCAGTGCAAAAGGCATCCTCCAAGACAGGGATCAAGCAAAAAAGTTATCAACCATCTATTATCATTGCAGGTCCTCAAAATTCTGGAAAAACGAGCTTGCTTACGCTGCTAACCACAGATTCAGTAAGACCAACTGTTGTTTCTCAAGAACCGTTATCAGCAGCGGATTACGATGGTTCCGGCGTCACGTTAGTGGACTTCCCAGGCCATGTCAAGTTGCGTTATAAACTCTCAGATTATTTGAAAACAAGAGCCAAATTTGTTAAAGGGTTGATAT tpg|BK006944.2|:160395-162555 7X198= 498=7X 
 tpg|BK006944.2| 338229 + tpg|BK006944.2| 338725 - INS CTTATATATATATTGTTACTACTGGACATATGAGTTTTTCTTGTAGCTTCAAAAGATCAAATATAAAATACGAATGTTTCTGAAATTACTGTAAAAGACTTAGGAAAAGGAATGAAACGTTTATATGGGAGAGAACGAAAATTTTTCCTTTTCCCGCCACTACTTTTTGCCACCATTTCCCGTTATTTATTTGGGCGAGTGCTCACCTCCGACGGAATCACGGG tpg|BK006944.2|:337767-339187 7X13=205S 10S193=7X 
 tpg|BK006944.2| 334247 + tpg|BK006944.2| 334793 - INS ACATTAACCAGTAATTGCTGTTCCACTTCTTGTATCGTTAAAGTGTATCTCTGATTCATAGAAGCATTTGGTAAGTGTATATTAATTGTCTTCCCATGGTATGCGTCACTCAAAGGATAAAATGTCAACAATGTTGATCTTGAGGAAAAATGGTAACAGATATACTCAGAGTTACTCAATAACAAACAATTGG tpg|BK006944.2|:333847-335193 7X10=86S 91S6=7X 
 tpg|BK006944.2| 299531 + tpg|BK006944.2| 299430 - INS GTTCAACATAGGGTTATGTTGCTCTTCCCGAAGATCCTGAGGAATGGCCATGTTGTTTGAAGAAATACCATGAAGAATTGTTGAAGTTTTCTAGTCCAAAAAAGACTGCCAAAGGAACTTTATTTGTTACAAACCTTTCTTCTTTCAAATCTACGCTAAACTTATTGCATGTTGAGTGTGGTAATCTAAAGAAAATCTGGAAAAACTTCAAAACCAACTACGACCTAAAGAGATTACATTGTGGTGGTCGTTCAGCTCAGCTGTTAAAAAAGACACCTAGTGCCTCAATAGCGAAGTTTGCACAGTTATATAA tpg|BK006944.2|:298790-300171 7X173= 294=7X 
 tpg|BK006944.2| 57783 + tpg|BK006944.2| 57727 - INS CCCTCATGCCATTATCAAACTCATTAATATCAGTTACCGAGGAAGCATCACTTCCTTCCTGTTTCTTTTTAGAGACAGATGTTAGCATAGAAATGACTTCAAAATTGGCCAGTGCCCAGTTATGCCACGCTTTGTACCATGTGTTGTCAAAATGTGTAGCGAGCAAATAGGAGCCTAGGATCGAATCTGGATTGCTCAATCTCCATTTAGGCTGTAAGCAAACTCTCCATTCTCCTTGCTTCAAGAAACAACGAGCTAAAAGCTTAGTATAATCTTCAACGTGACGAGGGACTCTTTTGCTTTGTTGAGGAACGCTTTGAGCTATCATATTATTTGGATCCAAACCTAAATCATGAGCCATTCTAGATGTGAAATTAATTAATTGCTTCAAACCCTCATCTTGCAACCCCGTAGCCCACAAGTACTTCAGTTGTGCAT tpg|BK006944.2|:56837-58673 7X154=1X343= 173=1X45=7X 
 tpg|BK006944.2| 360615 + tpg|BK006944.2| 360490 - INS TTTCTTGCTCATTGGTTAGACTACCTCAATTGAGAAATACGATGATTGAATTAGAAAAGGAACTTATGAAATCTGGGATTATAAGTGAAATGGTGGATGATACCATGGAGAGTGTTGGGGACGTAGGGGAAGAGATGGACGAAGCTGTTGATGAAGAAGTTAATAAGATAGTTGAACAATACACAAACGAGAAATTC tpg|BK006944.2|:360082-361023 7X5=192S 185=7X 
 tpg|BK006949.2| 528473 + tpg|BK006949.2| 528338 - INS GTATACAACGTAGCAATATCATATCGTCCCCCTTAGCTAGTACTCGTTTACCTACAGCAAACGTGTCCACTGAAGAATCCTCTATTTTACCAAATGAATCATTGAAGCTAAAAAGAGATTTATTGCGTCTTAAAAGGTAAATAGTGCCGAACAGTCAGGAGCACACAATACATGACCTATAATGACACTATCTTAATG tpg|BK006949.2|:527928-528883 84S262= 99=7X 
 tpg|BK006944.2| 30451 + tpg|BK006944.2| 30918 - INS GCATTGTTTCATTCTTCGACAGAAGTAGGAGTGTTATTCTTCTCACGGCCCTTGTTCTTTTTGGAGACTCTGTTAGGCTTTTGGCGATAATGGCTCCCTGGCCTGCCTCTTCCGTGTTCTTGAGCCGTCTGTTTGCGACGGTTGTGGGCATTCATTCTAGAATGCTTTCTCTGT tpg|BK006944.2|:30089-31280 7X7=14S 153=7S 
 tpg|BK006949.2| 339453 + tpg|BK006949.2| 339655 - INS CCATTCAGCGGCGGTCAGGGTAAGCTTGGTGTCGAGAAGGGCCCTAAATACATGCTTAAGCATGGTCTGCAAACAAGCATAGAGGATTTGGGCTGGTCTACGGAATTAGAGCCCTCAATGGACGAGGCCCAATTTGTGGGAAAGTTGAAAATGGAGAAGGACTCCACAACTGGGGGTTCCTCTGTTATGATAGACGGTGTCAA tpg|BK006949.2|:339033-340075 7X72=29S 3S1=444S 
 tpg|BK006949.2| 874069 + tpg|BK006949.2| 874412 - INS GGGTGTATGGCTTTGTATGATGTTTTACATGGTGAGAGGCACGTAAATCGTTACAGCGAAGGCATACGGTCGGAGAATGACGAAGCAGAGGTTGCCCTAAGGCAGCGTAGAAATTTACTACTCTTTTGGCGAAACCACTCTTCTACACCAAAACCTTCACTACGCCGAGCCGCCACTATAGTATATGAGGATCATGTATCATCCCGTTATTTTGAGGATATAAGTTCTATATTAGGAAGCACTGCAATGAGAACTAAAAGACTATCTCCCTATAATGCGGTAGCATTGGACAAGCCTATTCAAGATATTAGTTACGATCCCGCAGTACAAACTTTATATG tpg|BK006949.2|:873375-875106 7X161= 170=7X 
 tpg|BK006944.2| 506517 + tpg|BK006944.2| 506806 - INS AAAATATTCAAGAGAAAGAAGAGACTGCTTACAACTGGTGGTGGTTCATTACCTACGAATAATCCGAAGGTTTCTATTCTGGAAAAGTTTATGGTGAGCGGGTCCATTAAGCCACTGTTAAAACCAAAGGAAACCGTTCCCAACACAAAGGAGTGCTCCACGC tpg|BK006944.2|:506177-507146 7X4=77S 78S4=7X 
 tpg|BK006949.2| 525033 + tpg|BK006949.2| 525676 - INS CCCATTGATAATCAAATTGCCGCGCATGCTAGATGAATAAGGAAAAAAAAAGGGGGACGGAAAACATTGCAACCAACACATTATTCTTTAGCGGCTTTTTGTGAAGAAGAGGAGTTGCTTGCTCCATCTTCATCGCTGTCATGGCCATTGAGACGCTGTAGCTTCTTATCCTTCTTGTCTGCACTCTCATGTTCAGATTGATCCAAACTCAAATTCTCTAAATCATGTACAATTTCAAGTAATTGCTCTTTAGAGT tpg|BK006949.2|:524507-526202 7X4=203S 240=7X 
 tpg|BK006949.2| 112200 + tpg|BK006949.2| 112345 - INS CGTCCATACACGAAATGTACAAATACGTACATGTTTCTGAGGTTGGTAACTGTTCTGGTTCTGGTATGGGTGGTGTTTCTGCCTTACGTGGTATGTTTAAGGACCGTTTCAAGGATGAGCCTGTCCAAAATGATATTTTACAAGAATCATTTATCAACACCATGTCCGCTTGGGTTAATATGTTGTTGATTTCCTCATCTGGTCCAATCAAGACACCTGTTGGTGCCTGTGCCACATCCGTGGAATCTGTTGACATTGGTGTAGAAACCATCTTGTCTGGTAAGGCTAGAATCTGTATTGTCGGTGGTTACGATGATTTCCAAGAAGAAGGCTCCTTTGAGTTCGGTAACATGAAGGCCACTTCCAACACTTTGGAAGAATTTGAACATGGTCGTACCCCAGCGGAAATGTCCAGACC tpg|BK006949.2|:111350-113195 7X330= 405=7X 
 tpg|BK006949.2| 546826 + tpg|BK006949.2| 546865 - INS CTGTTATGTTAACGCAAAAGAGGCTCATAATCATTATCTTCTCGGCTTGGTTTTTCACATCTCTGGTTTTCTTACCAGAAATTCAATTTGGGCTAGATCAAACATTGGCTGTTCCACAGGATTCCTACCTGGTTGACTATTTTAAGGATGTTTATAGCTTCCTAAACGTAGGACCACCGGTTTACATGGTCGTGAAGAATTTAGATTTGACTAAAAGACAAAACCAACAGAAAATATGTGGTAAATTTACAACTTGCGAAAGAGACT tpg|BK006949.2|:546278-547413 7X3=212S 134=7X 
 tpg|BK006949.2| 200217 + tpg|BK006949.2| 200433 - INS CGATGGGAACCACCACAAACTTCACTAGCTAGTTCATAACAGTTGGTTTCATTGTAGAGATAAAACAAGCTGGACTTGAACCCATAAGTAATGTATTCACCTTTTGAATTAAAGAAAGCGCCCTCCAAGAAACCTTTCATCATCTTATTAGAATGCAAGACCTTATAACTTAGTCGGTAGGGACCCTCTTCCAAACTGTTTTTCGTCAACTCAATAAATACATAATAGCCATCCCTATTTGTTACTGAGAAG tpg|BK006949.2|:199699-200951 7X126= 275S3=7X 
 tpg|BK006944.2| 611870 + tpg|BK006944.2| 612585 - INS TCATCTCATATACTCCCAAGCTTCGAAATTAATCTTCGATCTATCTACTCTGGAAAAATGCTTTCTTTGGCCCTCTTTGATCTCGTCGGTTCCAGCAGGAATGTTCAATTTATTGGCGCTTGATGAACTGGAAGCAGATGGAGTTGATTCGTTAGATGAGGCAGGCGTTTCTTCGGCCTTGGATTCGTCTGCAGTTGCTTCTTTTGTTTCCAATTCAGAGCTAGAACCAGAGTCTGAGTCGGAATCCGAATCGGAGGAATCAGAAGATGTGGATTCGTCGGAACTTGAATCAGACGAGCTTGAAGAATCGGACGAGCCTGAAGAGTCTGAGTCCGAGCTTGAGTCGGAATCCGAATCTGAATCCGAGGAAGAGCTGCTAGAGCTGGAGCTAGAGTCGGAGTCAGATGAAGAGTCGCTGGAGCTGGAGTCGGAGTCAGACGAAGAGTCGCTAGAGCTGGAGCTAGAAC tpg|BK006944.2|:610922-613533 7X161= 256=1X196=7X 
 tpg|BK006944.2| 414055 + tpg|BK006944.2| 414625 - INS TTTCAAAGTTATACTCTTTTGCCATATCGACGTACTTGTATGGTGTTTTTACGACACGAGATATAGTTTCGTCAAACCACTTCCAGACTTGTTCCATGTTGTCAATTTCAGAAACTTGAAGGGAAAGCCCTTGAAGACTATTCACTAAAGCCATCACTGGTGAAATTAAAGATATGTTGAAGATAACGTTTGTTCTCGTCAGCTCATCGAGCAAGTTGGATATTCTTGTAGTTATCACGTTAGAAGCATTTTTGGAGGATGCTAGCTTTAATAGTAGGGTGAATAAAGAATTTCCACCAGAACTTGGATTCCACCACCTGGTTTGAGTAGAGTTAAATTCTTGAAATTGTAAGTAGTTGTCCAGAAT tpg|BK006944.2|:413307-415373 7X230= 184=7X 
 tpg|BK006944.2| 540329 + tpg|BK006944.2| 540537 - INS CCTTAAGAATATAATACCCCTTTTTGAATTGAGCAAGTCATAAAAAATTTTCTCATGCTTAATCGTATCAATTGTAGGAATAACAATGTCAGGCCTCATGACCTCATGTGCTTCTAAAGAAACAGAGGGAATTTCGGAACAAAAGGAACTAAAACTCAACTTATCGTTCGCAATAACTATGGTAGAATAATCTGATAGTTCTTGGCTGTCATGTCCAAAATAAGTGTTTATAGTTTGTATAAAAGCTCTTTGTGATTCACCAGTTGAATCACCAGCTAGTGCATATAGTAGGGATCTCTTAATC tpg|BK006944.2|:539707-541159 7X218= 285=7X 
 tpg|BK006944.2| 386539 + tpg|BK006944.2| 386077 - INS TTCAAGATAAATTAAATAGGTTAATGGACCAAATTCAGCCAATCATTGATTCTTTGAAAAAGATTGATGATTCAAGAATTGAGGAGAATACTTTCGAAATTGCATTGGCTCGCTTGATACCACCTCAAAATCAATCACATGCAGCATACACGTACAATCCAAAGAAAGGCAGCACCATGTTCAGACCGGGAGATTCTGCTCCATTGCCAAATCTTATGGGTACTGCTCTTGGTAACGACAGTAGTAGACGTGCCGGTGCTAACTCTCAAGCCACATTACACATCAACATTACCACGGCAAGTGATGAAGTGGCTCAAAGGGAATTGCAAGAGAGACAGGCTGAAG tpg|BK006944.2|:385373-387243 7X212= 173=7X 
 tpg|BK006944.2| 34772 + tpg|BK006944.2| 35138 - INS ACACCTTACTATCACACATGAATATATATATATAAAATAAGCCAAGACAGTGGCCTTCCCTTATTATCAGCGTACTAAAATCTCATATGATTTATTTTTCGTGGTCCTGAACGAGTGTGAAAAATTTTGAAAAACTCGCAAAGGAAATGCCAAGGTCAGCAACTTT tpg|BK006944.2|:34426-35484 47S13=30S 77S6=7X 
 tpg|BK006944.2| 372794 + tpg|BK006944.2| 373207 - INS AGAAAGAGCAAGATCTAGCATTGGAGGAAATAGAAGTCAAAACAAAATGCCATTATTGTGGAGTTTTGTAATTGGTACAACAATAATTAGAAGCTTGCCCGTTGTGTATGTTTTCACTTACTCCTCTAATGTGTTCAGGCACCATAAAGATGTTCATTTCGTCGTATTTTTATCATTGTGGCTACTGTTTCAAATTAGTATACTGTATTCTCAAGATGTATTGGGATCGCGCTGGTTCTTGCCTAAGCACACAATACCTGATGGATATTCGTATTTCAAGCCCCTTTCAAACGAGTATATATCGG tpg|BK006944.2|:372170-373831 7X249=17S 1S1=230S 
 tpg|BK006944.2| 293282 + tpg|BK006944.2| 293282 - INS TTCCTCGAGAGGGCTGTTTTTATCTTCCGTCACACTAATAGAAAACCACTCTATCCAGTTTTTTTTGTTACTTAACTTATCTTAACTCGATATTGTATAAATACTGAAGTCCATATACTTCTTTTTTTCTCCTTTGGATAGTAAATACGGTAAATTAAAATTAGTGTAAACTGAACAATATTAACATAT tpg|BK006944.2|:292890-293674 7X5=89S 89S6=7X 
 tpg|BK006944.2| 276075 + tpg|BK006944.2| 276268 - INS ATATGGGCCAATGGTATATGTAACAATTTGCTAACTTCTGTGATGAGAGATTGGTCACCACTGACCCCAGTGTTGATTGCGCCTGCAATGAATACATTCATGTATATCAATCCTATGACAAAGAAACACCTGACGAGTTTAGTGCAAGACTATCCGTTCATCCAAGTTTTGAAACCGGTGGAAAAGGTATTAATATGCGGAGATATTGGTATGGGTGGTATGAG tpg|BK006944.2|:275613-276730 12S205= 4S6=1X3=7X 
 tpg|BK006949.2| 451159 + tpg|BK006949.2| 451644 - INS TTGAAGATTTTAGTAACACTATGTTTGTATTGGAATCTTTCCTCAATCGTTTCTGCTGCCTTGCCAGCAAAGTGGCACTGGCAGTATCACTGGTACTTTTACTCAACTTTAGTCTTAAGCCTAATGAATTTAGAATTGTGACAAATCTTACTTTTATAGCATTAAGTTTCCAATTTTTGGTTAGATTACTGAAATTCTTGGAAC tpg|BK006949.2|:450737-452066 7X87=15S 1S1=258S 
 tpg|BK006944.2| 91488 + tpg|BK006944.2| 92104 - INS CTTTTAATAAGTCCAGAACCAAAGTAGTTGAGTCACTGGAAGAGTTAGAGCTTGCGGAAGACAGCGAAGCAGAAACTAACCTTGAGAGGCCATCTAGTGTTTCAGTTGCGTTGTCTGAATACTTCAGCAGCCCATTAATCTCTGTCAACTGCCTCGTGCTA tpg|BK006944.2|:91152-92440 7X5=75S 76S5=7X 
 tpg|BK006944.2| 412901 + tpg|BK006944.2| 412474 - INS GTCAATGTTCGTAACTTATATTGGCAACGGTATGACAATCGCTTAATGAGCAAATAATAAACTGAAATATTTTGCAATCAAGGAAATTTTCAAATTCATATCTGTATGTTACATTGCCCTCGTCATCTTTGACCATTTTTACCAGCTCTTTGTTATGGATTATTAATAGCAGTAAAAATAATGGATCGTACATATCAACACCAGATCGTTCGGTATCATCGTAGTACTTTTTGACTAGGTCACACC tpg|BK006944.2|:411968-413407 15S13=174S 123=7X 
 tpg|BK006949.2| 218503 + tpg|BK006949.2| 218444 - INS CTCCTATTTCATAAAACAATGGGCTTCAATATAGCGTATGTCTAGCTCACAGCATGTGTTCCAAATACATTAAAGAAGATCTCTTTTGTGGTTGATACTAACCAGTAAAGTTGAGAGTTATAACAATGAAAATAGGATGCTGTGCGACTTTTTTTATCCACAGTTAGGTGGAGTCGAATTCCATATATATCATTTATCGCAGAAACTAATCGATTTGGGCCATTCTGTCGTCATTATAACTCACGCTTACAAAGATCGAGTCGGCGTACGACATCTTACCAACGGTCTAAAGGTCTATCACGTACCATTTTTTGTGATTTTCAGAGAAACCACTTTCCCCACTGTTTTTTCAACATTTCCAATAATAAGG tpg|BK006949.2|:217690-219257 7X262= 78=1X280=7X 
 tpg|BK006944.2| 154718 + tpg|BK006944.2| 155031 - INS CCTAAGAAGGTTCTTCTCTAATAGGCAAAGCTCACCCTTGTTTAAGGTCTATTGCTGCACACCCTAGGTATTTATCTAATGTGTACTCACCACCAGCAGGCGTCAGTAGATCACTGCGCATCAATGTAATGTGGAAGCAGAGTAAATTAACTCCCCCAAGATTTGTGAAGATCATGAATAGACGCCCTCTGTTCACAGAAACTAGTCA tpg|BK006944.2|:154288-155461 7X153= 104=7X 
 tpg|BK006949.2| 361944 + tpg|BK006949.2| 362011 - INS ACTATCGATCTTTGGGAAGATCATTATAAGAGGTCCCAAGCCAATTCGTTCTCAAATGCGTCAAATACTGGTACTTTGGAGGGAGATTCTGCAAATTTGAACAGGGTGGCTACCAATTTACTAGCAAATGCCACTCAAAAAAGTGTGAATGGATCTAATCC tpg|BK006949.2|:361608-362347 7X5=75S 77S4=7X 
 tpg|BK006944.2| 308644 + tpg|BK006944.2| 309357 - INS GATCCTTACTCCTTGTTATAGTATTTTTCTACCTGTTGATTGCAAGTAAGGGCAGCATTATCCTGATAGGAGTAGAGGTTAACCGCACATCGGAATGAGACTTCTCCAAGAACGTTCTCAAAGTAAAACATTTAGCATTAGGAAATTTCTTTGGTCGATTATTAGACAAAGATTAGAGTGTATTATGTTCTGATGCTTAGTTAGAACGGAAAGTGTTACCCATCTTGCAA tpg|BK006944.2|:308170-309831 25S19=1X36=41S 109S6=7X 
 tpg|BK006944.2| 54539 + tpg|BK006944.2| 54816 - INS AAGGAAGACAGGCAATTAAGGCAAAATAAAAATCCAAACGGAACAAGAAATAGCAAGGGAAAACAAGAGGAAACAGCAACGCCAGATCTGCCTCAACAGCAATACATGCCACCACCCCCACCTCCAGGGTTTTTTCCAATGCATCCTAACTTTCCTAACGGCCCAATGCCACCATTACCACAGGGGTTCCCAATCCCACCAAATGGTATGTTACCGGTAACAGGACAAC tpg|BK006944.2|:54067-55288 7X88=26S 1S1=337S 
 tpg|BK006944.2| 633034 + tpg|BK006944.2| 633292 - INS TTTAGAATCAGTAATTCTACAATTAGGACAATCCCAAGCATTGTCGCCTGACAGTTCTTCATCGCCTGTAAATAAGTTTATGCAATCCTCTAATTTAATTTTTCTCGACTTACTTGTAAAGCTATACAATGATAGTTTTGGAATCGCAAGTGACAGAACATAGAAGGTAGAATAGCTATAAGAAGAATTACCACAGCGCTGACATTTCAAAATGTTCTCCAACGGCCCTCGATATATGTG tpg|BK006944.2|:632540-633786 7X194=16S 8S1=192S 
 tpg|BK006944.2| 8753 + tpg|BK006944.2| 9051 - INS GATATCATGCATCGAATCTATTATCTTCCAACCGAACTTTTACAAACGTTTAGACCGAGCGTTATTGACTGAATTAAGAGCAAGTTTTTACACGTGTGACTCTGGCACATTAGAGCTGTTTGAGAATCTAAAGTCTTGCTGTCTAAGGACCAAAAATAATGTATTTCGAGGTCATAGCTAAGAATCTCATTGTTCTT tpg|BK006944.2|:8345-9459 7X5=93S 94S5=7X 
 tpg|BK006949.2| 39083 + tpg|BK006949.2| 38795 - INS TATCTAAATAATGTACACAGTTAGCGTCTAATAATTAATTAACGATACCAATTTAATTCATTCACGTATTCCTCACCTCGTGTGTAAATTACTAACAGAGTAGTAATAATAATAAGAATCAATAATAATAATAAATCCATCCTTGTGTATTACCCGGGTTAGAGG tpg|BK006949.2|:38451-39427 7X5=148S 83=7X 
 tpg|BK006944.2| 96958 + tpg|BK006944.2| 97527 - INS GTGCAGATATTTTCGCCCATTTCGAAGTGAAATCATTCTAATAACTTCTCCTGCGCAATAGATTGGTCATCCTGATTTTTATTCTGAAATCGAAAATGAAAAGCATTTATTGCACTGAAATAGCGGAACCTGCTTCTAATAAGCTTAAAATTCAATCATAATAGTGTAGTTAATAGAAAGGACAGAAGAACTTTTCGTTCCTTGGTTTATCATCCAGGTTTCAGCACGGCTTTTGTTTCAAGTTTAAGTAGGTA tpg|BK006944.2|:96436-98049 7X3=288S 127=7X 
 tpg|BK006944.2| 281029 + tpg|BK006944.2| 281033 - INS ATCTTATTCTTCCTTCCTCCCTTCTTTTTACCTGTTTTTAATCTACCCTCAAATCCGGCTCTTTTCTTTGGTACGGCACTACCGACATACTTTCTTTTCATCTTTTCTTGCTTATTTCTCTTTTTACCCTTGTTGTCTTTCCTAATCCTCAGATTCTCTTCTCTTCTCTTTTGTCTTTCAGATATCGTGTCTTCCACAACCCTCTTACGTT tpg|BK006944.2|:280593-281469 7X177= 185=7X 
 tpg|BK006944.2| 259985 + tpg|BK006944.2| 260694 - INS GATGCTGAGATCTTATACGTTTCTTTCTTTCGCTATCTTCCTTGAATTTTTTTTCTGTCTGAAGTAAAATATCCCGTAACAAACTAATAAATACTACGAAAGTCTCAAAAAACAATAATGAAATTCTCCACTGCTTTGTCTGTCGCTTTATTCGCCTTGGCTAAGATGCTCATTGCCGATTCCGAAGAATTCGGCCTGGTGAGTATCCGTTCCGGCTCGGATTTACAATACTTGAGTGTTTACAGT tpg|BK006944.2|:259479-261200 15S7=1I107= 45=1X17=67S 
 tpg|BK006944.2| 504372 + tpg|BK006944.2| 504422 - INS CTCGTGGTCCAAAGAGGTAGACCTTATGGTGTGTTTTGAAGATAATTGAACTCATCCATTGCTTTAACGAACTCTCTGATTTGCAAATAATTTTCAGTTTCCTTTCACTGTTTTCTAGGGTCAATAATAATAGTTTTGAAGATATATTGGACTTCTTTTGGTGTGTTTTCGATTTTCCATTCTTGTCTAGGATATTAT tpg|BK006944.2|:503962-504832 7X11=1X273= 16S158=7X 
 tpg|BK006944.2| 89419 + tpg|BK006944.2| 89184 - INS TTAAACACAACACCATATTTATCATCTGCCGTACCGCTCTTTATAATGGCAATCATAACGGATATGATAATGGCTGCCAATACAGTGGCTACACCAACGCAAACGTGTAGAGCTAGGGCAATGAGCCATAATGGTTGTTTGAACATATATCTGT tpg|BK006944.2|:88862-89741 7X64=51S 1S1=175S 
 tpg|BK006944.2| 622609 + tpg|BK006944.2| 623334 - INS CATATTGGAGAAACATGAACAATTGAGCTCAAGCGATTATGAGAAGCTAGAAAGCGAGATAGAAAATTTGAAGGAGGAACTAGAAAATAAGGAGCGTCAAGGAGCGGAAGCCGAGGAAAAATTTAACAGGCTGAGAAGACAAGCGCAAGAGAGATTAAAAACATCAAAACTCTCACAGGACTCATTGACTGAACAAGTAAATAGTCTAAGGGATGCAAAGAACGTGTTGGAAAATTCCTTGAGTGAGGCAAACGCGAGAATCGAAGAGTTACAAAATGCAAAAGTAGCACAAGGTAACAACCAGTTAGAAGC tpg|BK006944.2|:621971-623972 7X156= 224S3=7X 
 tpg|BK006944.2| 620372 + tpg|BK006944.2| 620617 - INS ACACTGACGAAGCAGATGAAGATAATGAAAATTTATCTGCAAAATCTAGTTCTGATTTTATATTCCTGAAGAAACAATTAATTAAAGAAAGGCGTACCAAGGAACATCTTCAAAATCAAATTGAAACATTCATCGTAGAGTTGGAACATAAAGTGCCCATTATAAACTCTTTCAAAGAAAGAACTGACATGTTGGAAAACGAATTGAATAACGCTGCATTGTTACTAGAGCATACAT tpg|BK006944.2|:619884-621105 7X1=1I200=16S 1=190S 
 tpg|BK006944.2| 397929 + tpg|BK006944.2| 397925 - INS GTCGTATTCATAAATAAGCACCCTATCCCTTAAACCCACGGCAAAATAATCACCTTTGGCGCCTAACCATCTAACACAAGTCCCGTTTGTATTATATTTTCTTAGTTTTAGTACAGCAGCATTTCTTAGAGTCATCAAATTCCAAAGACGTATAGAATGGTCATCACTAACACTGATGGCAATTCTATTGGTGGGGTGAATATCCACATCATTAACCCTTGCCGTGTGTCCCTTTAAAGTCCCCACTGTTTCCCAGTCCTTTACTCTCCAAACCATAATTTTGTGGTCTTCTGATGCTGATAATAACCATTTGCTATTCTTGCTCCCCTTTGAAACAGCAGCATCCTCACTGGAAGAAGCTGGATGTGAGAATTGTAGAGCAGTAATAG tpg|BK006944.2|:397133-398721 7X170= 195=7X 
 tpg|BK006944.2| 196409 + tpg|BK006944.2| 196995 - INS GTCGTATGCAGGGTTTTGAGCTGTGTTTCGAGCTTACTTTTGCAGCAGGGATTGCAGATGACTTTATTGGTACGGTCTTATCCGGTTTAGGATTGTATGCTGCCTGTGCAGCGGTAGCTGCCAAAGATAACGGATTCACAGGTTTTTGCGAAGGGAGAGGTTGCTTTTTTGCAGCATCCCTATGACTTCTATGGCTATGTGTATGCTTATGAGTAGATTTGTGTTTACTCTTTTTGCTTTTGATAGGTTTCCCGCTCAACCCACCTGGATTCTTAGGTTTTTTATTCGATTTGGAGTTAGCAGGGTGTCCAC tpg|BK006944.2|:195771-197633 7X5=72S 293=7X 
 tpg|BK006949.2| 66600 + tpg|BK006949.2| 66791 - INS ACGAATTTCGTGTACTTCCGTTGAGACAAATTTCGCGATGATTTCCGTTTTCGGAAAGATGGAGCCGGGTAAAGCGCGCATGAATTGATAACTTGGCACTTTTGAACCTCAGTATCATTATTAACAATGTATAGTTGCTTTAGTTCGCATTTCAGGGTAAAAGTGCGGAGGATACGAAAAAGATGAGATAACTTACAGAAGGAAACGAATAGTGGTTTCAAAAAATGCCTTTCACTCGTAGAGAAAACAATAAAAGTTACCGCACTCCAACACAGGCGATACTGGAGGAATATTTTCAAGAGTAAATAGAAGCAAAGATGCTTAAAAATGGATACTTGAACCAATTTTTCTGTAGCGGTATATTAC tpg|BK006949.2|:65854-67537 7X354= 12S1=216S 
 tpg|BK006944.2| 355630 + tpg|BK006944.2| 355764 - INS CTGTAATGCTGTAGAGCGTGCGTGCGATATTATTGATGGATATCGTCTTTATCTTTCCGTGGACCTAAAACGGCACCCCTTCGTCTAGGATAAACGCGGTCGGCTCTTTCGAAGACTAAAAAAGCAGCCACAATAACGTTACATGCAAAATCAGCCCACTCGAAGTTAGATACTGCGTAGACGGATTTGCACGATGCGATGATAAATATTAGGGACAGTGCGTGCCCACCCATAAGTTGCTGTAGAGCTTACAAATTGTAAAGACTAATTCCAATCGCACGCCCACCCCTCACGGGAATAAGTTAGAATGTTGCGGAATGAACGATAACTTCATATTAGGTAAAAGGGAAGAATGCAACGCTGCGGTCTACGGGCTTTTTTCTGCGAGACCAATTTTCTTCTTTTGTTTTTTTATTTCGATATTTAGTTTTCATGCAAACGGGTATTATTCTTGACAGGCCATTATGTAAGAGTGTGGAAACATAATTCTTGCACATACGACGTTTTCTTAACTGTTCCTGTTTCAAGTTACGGAAACGCCTGTGGCCCAGGTAGCGTAGGCAAAATCAAGCTCAGAAT tpg|BK006944.2|:354458-356936 7X160= 2S559=7X 
 tpg|BK006944.2| 43726 + tpg|BK006944.2| 43806 - INS TAGAGTCATTTCTAAGATCCATAACCCAGTATTCACTGCAGCAATCTAATAGGAATCCTTTAGCAAAATTGAAAATACCATCTGCCGCAGCCACACCAAGAACAAGAAGCGACCATTTCGCCAAATAATGTGAAGAGCCAGTTTTTCCATCCGTGGATGGGACAATTCCTTCTAGTAAGAAACTGAATGTGTATGAAAAGACGGGATTTGTGGCGC tpg|BK006944.2|:43280-44252 7X286= 108=7X 
 tpg|BK006949.2| 505960 + tpg|BK006949.2| 506701 - INS AACCGTGATAAACACTCCAATCATTGTGGCCAATTTATTGCATGTTTTAGCTACACCAACATCCATTAACGGACAACTAAAGCGAGCGCTCGTCCTAGTGTTGAATGCAAAACCTATAGATAATGTAAGAATCAAGGAGGCCTTAGAAGAGCTGTCGTGGTTCTCTAATACTGGGAAGGACGACGACGATACTGCTGTCGAGAGCGATGATGAACTTTTTGAAAGGCCTTTTAACGTAGTTACCGCGGACTCGCTGAGCATTGAAAAGAGAAGAAAGCTATATATTTC tpg|BK006949.2|:505370-507291 29S122= 113=38S 
 tpg|BK006944.2| 11812 + tpg|BK006944.2| 12540 - INS GCTCCAGTTAGGAAACCTTAAAAAAATATGCAAGGATTCTAGATTTCAGGCTAGTCTTCAACCACTTTGCACTTCCGGATTAAAGGCTTTTATAGAAAACATCTTGGTTTGGGACTATATTGCTAGGTGAAAATTTCAAAATTGTACAAAAGATCATTCTTGTTTTTTTGCCTCATTAGCTGATACAATGCGGAACTACATGGCGCTCTTTTATAAGCATCTACT tpg|BK006944.2|:11348-13004 7X333= 211=7X 
 tpg|BK006944.2| 424259 + tpg|BK006944.2| 424470 - INS TCGCTATTCTTTCGATTAAATCCAACGAAAACAAAGTCTCAAATTTGTCAACCCCATGCAACGCCCCGCAAATACCGTACATGGCATTTACAAGCCTGGTTAATATTGGTTGGTCTGTCGCATTCGAGAAAATTGGCTTCAGCGTTGGAAGTACTTCAACAATGGTCTTAAAGTCATCCGTTCGGATACTGCTACAGGCGTTCGAAACAATTGCGATAGCCTTCCTCTGCGCATGTA tpg|BK006944.2|:423771-424958 7X8=8S 119=7X 
 tpg|BK006944.2| 329867 + tpg|BK006944.2| 329858 - INS ACCGCTTATACACATTTGACAAAGTGGTGGCTGAGACTTTAAAAGACAATACCCAATCTAAATTGACTGTGAAAGGAAACCTGGACACATATGGATTTTGCGATGATGTTTGGACTTTTATCGTAAAAAATTGTCAGGTTACTGTTGAGGACAGCCACCGCGACGCCTCCCAGAACGGGTCTGGAGATAGCCAAAGTGTAATTTCGGTGGATAAGTTGAGGATTGTGGCATGTAACTCAAAAA tpg|BK006944.2|:329358-330367 18S76=34S 117S5=7X 
 tpg|BK006949.2| 769054 + tpg|BK006949.2| 768322 - INS AACATTCATATGGAACGGCTTTAGGTGTTATCCGTTCTTTGTGGAAGGATTCACTTGCTAAAACCGACAAGGCAGACTCGGGATTGGACAATGAAAAATGCCCGAGGATGGGCCATGTCTTCCCACTGGAAACTAGACCTTATAATCAAGGGTCAAGGCTAACAGCATACGAGCTAGTTTATGATAAGATTCCATCAACTTTAATTACTGATAGTTCCATCGCGTATAGAATTAGAACTAGTCCAATTCCAATCAAAGCAGCATTTGTTGGAGCTGATAGAATTGTTCGTAATGGGGATACAGCAAATAAAATTGGTACTTTACAACTTGCTGTAATTTGTAAGCAGTTCGGAATTAAGTTTTTTGTAGTAGCTCCCAAAACAACTATCGATAATGTAACCGAAACTGGCGATGACATTATTGTGGAAGAACGTAACCCTGAGGAATTCAAGGTTGTTACTGGTACAGTAATTAATCCTGAAAATGGTTCCTTGATATTGAATGAGTCAGGAGAGCCAATCACTGGAAAGGTCGGTATTGCCC tpg|BK006949.2|:767222-770154 7X4=161S 272=7X 
 tpg|BK006949.2| 747560 + tpg|BK006949.2| 747669 - INS GGGTGCTACTGAGAGGGACATACTAACCACAACTAGATCTGACTGGCTTGTGAAGTTGCTTTATGCATTTCAGGATCCAGAGAGCCTATATTTAGCAATGGAATTTGTACCGGGTGGTGATTTTCGCACATTGTTAATAAATACAAGGATATTGAAGAGCGGTCACGCAAGGTTCTATATCAGCGAAATGTTTTGTGCCGTGAACGCGTTGCATGAACTTGGTTACACTCACCGGGATTTAAAGCCGGAGAATTTCTTGATTGATGCTACAGGGCATATCAAGCTGACCGATTTTGGTC tpg|BK006949.2|:746948-748281 7X265= 150=7X 
 tpg|BK006949.2| 213066 + tpg|BK006949.2| 213511 - INS TAGTTGTCCAGATGAAGCATTGAATGCCTTAAAATATTTGTCCGATACAAAGTTAGACGAAAAGACAATTACCATTGATCTAGATCCTGGTTTTGAAGATGGAAGACAGTTTGGTCGTGGTAAGAGCGGTGGTCAAGTCAGCGATGAATTGAGGTTCGATTTTGATGCATCCAGAGGTGGCTTCGCCATTCCATT tpg|BK006949.2|:212662-213915 7X5=92S 94S4=7X 
 tpg|BK006944.2| 151039 + tpg|BK006944.2| 151501 - INS GGATTGAGTAAGATGTGGGCCTGAGTTTCCTGTTAGAAACAAAGATATGCTTAAAACTAAATAACATTGGAAATTAGGGCATAGTCTTCAATGTTATACTTAAACATCACAGCAGGAGATTGAGATGATTGAAAGAATGGTGCAAGAAATGATTCATTAACATTCTTCCAAGTTTTGCAATATTTGCAAGTATTACTATCAGACTTTAGTTGAAGTGACTATGCTATTACCAAATTTCACTGGAGCCAGAAAAATAAAGATCACTTAGAGACAAAGAAAAGTAACA tpg|BK006944.2|:150453-152087 7X182= 269=7X 
 tpg|BK006944.2| 158928 + tpg|BK006944.2| 159650 - INS GCTTGAGAACCATCCCATGAAGTAGCGAGAAGTTTACCCTTCTTTAACTCTATACTGAATTTGGGACGCTTGATGCTTTTTTGAAAATTGCAGAACTTTAAGTCTTTACCCTCTTTATGAGTATAAAAGTTAGGATTTCCAACCTGTAAGGGACATTTCCTTTGATGTGGACAAGGT tpg|BK006944.2|:158560-160018 7X6=82S 83S6=7X 
 tpg|BK006949.2| 225155 + tpg|BK006949.2| 225423 - INS GGTCTCTTAGATCGGTAGTAGCTTCGCTTCCACTTGAAGTTGATATATCATCTGTGCATCTTAGCGTTTTCATGGCAGTCGATTCAACCTTTTTATTGCAATTAGAGGTTCTATCACCATATCCAAAATTGGGAGTAAATTCTATCGGCGCAGTGTTTATATGTTGCTGTTTCCCGCCATGATTCCGACTAATATAACGAACTCCATTAAATCGAATTTTTATTTGAGTATCGTGCAGCTGTGTACCAATTTGTAAGTATAT tpg|BK006949.2|:224617-225961 7X407=1X44= 246=7X 
 tpg|BK006949.2| 251754 + tpg|BK006949.2| 251832 - INS GAACCTCTCATGTCACTCATTTGCGAGCGAAAAAAAGAAACGGTAGACAGAATAGGCGTTTGTTATCGTCGATGGTGAGAAAAGGCGATATCGCCATTAAGGTAAACAATTATTATGATTATGGTTCTTATGGTTGATACGTTGATTTATATTAATATTAATGAATGCAAACTTATGTTATTATATATTTTTAAATTTTCATACCGACAGGAAGAGTCAATGACCTCTTGACCACACCTGTTGGTAGCGATATAATGCTGTTTGAGTAGGCAGGATTTAGC tpg|BK006949.2|:251178-252408 7X193= 3S58=1X202=7X 
 tpg|BK006949.2| 205726 + tpg|BK006949.2| 206005 - INS CATATATCCTTACTGAGTAACTATAATTATGGTTCATCGAGGAAGGACTTTGAAGTCAGACACTGATGTAACATCTCTTAATGCGTCAACAGTATCACACCAGTCAAAGCCATTTAGACAGTTTTCGACTAGGTCGAGAGCAAAGAGTAACGCA tpg|BK006949.2|:205404-206327 7X5=72S 73S4=7X 
 tpg|BK006944.2| 185502 + tpg|BK006944.2| 185451 - INS TGTTATACCGAATATCTTCAAGTTATCTGGAACAACTTTCATATATTTGATAAGATGGAGCAAAACAAAGATCCGCAGATGATCTCGAAACATAGTTCTAGGCTACCTATATGGGTGCTAAGTCCTCGCGAAGAACAACAG tpg|BK006944.2|:185155-185798 7X10=60S 65S6=7X 
 tpg|BK006944.2| 244163 + tpg|BK006944.2| 244642 - INS GTTTAACCTCATTAGGATAGTGACAAGATTTACATAATAACCCGTATGAACCTTCTAGTTCTAAAAGAACTAGCTTGGTTAATTCGTGGAAATCTAAGTCATGCCCATTTTGTAAATTTGTATTGTATAAATGCAAATATAGTTTAGCAATACACTCGGTATCGGTATCACTTTCGAATTTATAACC tpg|BK006944.2|:243775-245030 147S90= 94=7X 
 tpg|BK006944.2| 393854 + tpg|BK006944.2| 394062 - INS ATTAACAAGAGCCAGAGGAACAAGGAGAAGGACCGAAAGCGGAGGGAAAGAAGAACGGCAAGGAGAAAAGATGAAAGAAAGCAGGAAAAAAAGCAGGAAAAAAAGCAGGATAATAAAACATCTCAATCTTTTCCTTCCTCAACTGACATGAATGGACAGCCTATAGAATTTTGAATGCATTCTAATGACATAACTA tpg|BK006944.2|:393448-394468 7X88=59S 4S1=327S 
 tpg|BK006949.2| 457414 + tpg|BK006949.2| 457885 - INS AATTTAATTTCAGCAAATTTAATATTAATTAACTCAGGATCACCATTCATAGAATCAGTTATGGCTTGACGAATCATTTCTTGCTTCATTCCGTCAAGCTCCCCCTGACTAATAAAAACCCAAGGATAAGCAAAATTTTTGTTAAACTTCACCTGCACTTCATCAATAGATTGTAAGATTTGGGTCATGGAATCCCTTTCAGTAATTAGTGAGACAAAGCACGCCTTTGGTGGTGATCCTCTATGATTGATATACGAT tpg|BK006949.2|:456884-458415 7X263= 129=7X 
 tpg|BK006949.2| 450724 + tpg|BK006949.2| 450868 - INS CATCAACACCGACTGCTGTTAGGTTTTTAAAGGCAATACCAGAATCACCAGGTTCAATTCCCTGTTCCAATTGACGAGACCTCAAATAATGTAATAGTGAGCGCAAATCAAAATCTAAGTCATTAATTTCAAAAGAGTCCATTTCCTTCTTTGT tpg|BK006949.2|:450402-451190 7X5=72S 72S5=7X 
 tpg|BK006944.2| 266464 + tpg|BK006944.2| 266563 - INS GCTCCATACTATATCCAAATCTCCAACTGTGTTA tpg|BK006944.2|:266382-266645 7X3=8S 1S16=7X 
 tpg|BK006944.2| 68103 + tpg|BK006944.2| 68257 - INS GGATTCTGGCTAGGTCGATGCACTACGCCGCGCTAGAACTATGGACCAAGCTGTTGACAATGTTCAGATGGTGATGCACTACCCTGTGCGGGGAGTGGCCACGGACGCGAGCGGAAGGTGCGGAAGGTGCGGAAGGTGCGGGAGTTGCGGGAGGTTCTTCGCTAAGCGTGAGGGTTGCTAGCTGGGGCGGCGGGGATTCCCTAAGTGTAAAT tpg|BK006944.2|:67665-68695 7X12=164S 169=1X16=7X 
 tpg|BK006944.2| 96467 + tpg|BK006944.2| 96939 - INS GTCCAGTGGCTCATCACCCACTCGTCACACCACAAGAGTGTGCGTGTCGTGTCATTCGAGTGATTCGCCCTGTTGGAGGCCATCGTGGTCGCCAAGAAAGCAAGATCAGCTATGTAACTCTTGTGGTCTTCGATATAAAAAAACACATACAAGATGTTT tpg|BK006944.2|:96135-97271 7X4=75S 75S5=7X 
 tpg|BK006944.2| 117098 + tpg|BK006944.2| 116393 - INS CTGATAGACGACTCGTTGTGTTTTAAAGAAGGGCTTGGTTGAAAGAACTGAGAAATTGTTGGCCTTTTGTTGAACCAAGAACCGTACGAACCAGGTTGGCTTGAGATAGAAGACGATAGATAATGCAATGAACTACTCCCACTTTTGAAGGAAGATGGCTGAATAACTTCCGCTAAAGACTCACTAGAAGACACAGATACTGAAGTGTTCGAGTTCCTCCGATTGGGTATTTGCCATCCTTTCCTCAAAGAATGGAAATTGGGTGATCCAATGCTGTTAGAGCTCACATTACTGTTGTTG tpg|BK006944.2|:115779-117712 7X5=190S 150=7X 
 tpg|BK006944.2| 229567 + tpg|BK006944.2| 229958 - INS GTCTTACCAAGTTTCACCTGTTCATCAAGTATTCTTCATTTCTTTTTCCATCGCGATGACGATGACAAAACGGCAAAAAGTCAAAGAAAAAGAAAAAAAAAGATTTTTTTTCCATCATATGCAGAGAGAATATGTCCAAGCCAAGCGCAGTGTGCATGTATGCTGTTTTTAGCATATCGGGTGTGCGAAAGGAATGACATAATGATTTGCAACTAATATTTCCTTATATAAATATGCTTCTGGATATGAGTCTCATGAAACAAGTTCAGTAATTGCTTGTTTTACCCTTACTTTTTTCTTGGTTATGACTTGTGTACATAATAAATTGCCTATTTTCCCAAATTGTGTCCTTTTTCCTTTCCGGTTGGTATGAGATATTTCTTTTCAAAAATCAAAAGAAAACAACAAAGGGTTGATATTATGTAATGCAATACCTAGAAT tpg|BK006944.2|:228671-230854 7X116= 221=7X 
 tpg|BK006949.2| 374594 + tpg|BK006949.2| 374772 - INS CTCAAAAGCTGCCTTCACGTTTCAATCCTGTCGTACTACAATAAAAAAGAGATTGAAAACGAGACAGGAAAAGTGAAGAGAGTTTATACCTTCCACAAAGGTTTTTGGGGGATGACTTTCCCGATGGGTACTATGTCTTTAGGAAACGAAGAGTTATATGTGCAGTATAACCAGTACGTTCCCTTATATGCATTTAGAGTCCTAGGAACCATATACGGCGGTGTTTGCGTTTGTTGGTCAATTCTATGCCTTTTATGCACATTGCATGAGTATTCTAAAAAGATGCTGCATGCTGCCCGTAAATCTTCATTATTTTCAGAGTCAGGTACGGAAAAGACGACAGTTTCTC tpg|BK006949.2|:373882-375484 7X159= 7S332=7X 
 tpg|BK006944.2| 382528 + tpg|BK006944.2| 382921 - INS GCGTTGGTCTAGCTAGACGCGCAGAAGCGTTGGTGATGGTGTCCAGGCCGGGTAGCAACCCAGGTCTCGAGTCGCCCTCTCTTAGTGGCGACAATTCGGCTAGTTGGTCCACTGCAGCGGAGATCATCTTGTCTGTGATGGTGGTGGCACGCGATAGTACGGCACCTAAACCGATACCTGGGAAAGAGTAACAATTGTTGTTCTC tpg|BK006944.2|:382104-383345 8X10= 15=1X177=7X 
 tpg|BK006949.2| 351302 + tpg|BK006949.2| 351494 - INS TGCTTGTAGGATTTTCTCTGATGTCAATCTTGTATTTAGTTTTGAACTCATCGGCGAAATGTTCTGTTATAGCCAAATCGAAGTCCCTACCACCAAAATGCTTGTCGCAGGCAGTTCCTAAGACTTTCAATTGACCCTTCTTGAAGGCCATGATAGAACAGGTGTAGGAAGAGTGACCAATATCAACAAAGGCAACAATTCTTGGCTTTTCTTCGCCTTCAGGCAAATCAGTCTTGAAGATACCGTAAGAAACACCGGCAGCAGTAACGTCGTTGACAATTCTAACAGGGTTCAAACCAGCAATTCTAGCAGCATCAGCAATGTTGTAACGTTGTTCTTCGGTGTACCAAGGTGGGACAGCAATACAAACATCGGTAA tpg|BK006949.2|:350532-352264 7X224=1X236= 367=7X 
 tpg|BK006944.2| 213898 + tpg|BK006944.2| 214226 - INS ATATTGGTGCAGTAGGAAGGAGCTGACTCCAAAGAAAAGAGCCAAACGAAACATTTGAACATACCAGGCGACAGGAGCCGACATTCCTCTATTGCAGATTCAAAAAGAAGCTCTTCTAGAT tpg|BK006944.2|:213642-214482 34S256= 13S93=7X 
 tpg|BK006944.2| 76416 + tpg|BK006944.2| 75682 - INS GGATATTCTTTGTACTGCACGCCACCCAATAAGAAAAAAAGGGAAAAGGAGCCGAATTTTGGTTTAAAAACATATAATGCTGAAATTGTGGAACACCAATTACCAACTGGAAGTAGGCTCGATCCAAAGAGTGTATATTATCAGTAAAATGCTTCGCAACTTAGTCGTCAGGAATGCGTGCAGAAACAGGCCGTCAATTCAAGTGGCAAGGGGGTTATGCCGACACCAAACAAGAC tpg|BK006944.2|:75196-76902 7X5=226S 2S220=7X 
 tpg|BK006944.2| 637869 + tpg|BK006944.2| 638313 - INS CCACAAACACAAAGGGCGTTTAGTAAATTATGCGGCGATGTATAAAAGAGAAAGCAGGCAAAAAGAAAATGAAAAATGAGACTATGAACTTTAAGAATTATGTCTTGACTAATTTTTTAAAACCCATCATCCATGAAGAGTTCTGTTTGTATTGTTTACGTTTGATGTTTGAAGTGAATTTAATAGAATTGTTCCTCTTTTTTTCTTCTTTTTTTAACTATAATATAATGTTTAGTATATCAACAGTACTATTT tpg|BK006944.2|:637347-638835 7X183=39S 4S1=270S 
 tpg|BK006944.2| 530547 + tpg|BK006944.2| 531140 - INS GGTAAGTTGGTTGAAATTTTTATGTTTCAAATTGATTATTTTTGCCTCTTATTGGCAGAGCATCATAATCCAGGGTCTAGTGGTTACTGGAAAGTTGGGTACGGGAAACCAAGATCGAACCTCTGGATATGTGTACAAGAATGGGCTCCTGTGTATAGAGATGGTGCCTTTCGCCATCTTGCATGCAGTAGCTTTCCCTTGGAACAAATACACAGCATTTAGCAT tpg|BK006944.2|:530083-531604 14S18=1X34=52S 108S5=7X 
 tpg|BK006944.2| 94405 + tpg|BK006944.2| 94403 - INS CTTTGGCTAACGAAATACTTGGAAAAAAATCAAATACTGCACCAGCATCGCCACATCATATGGATTACAATCCAATTTCCTCATTAACACCAGGCAATTCACCAGAATTCAACAAGGCAAGCTTATCTCAGATTAGTTTTACAAATCCATTGAACTATGGGTCTGGCTTAGGTTTTTCCTCTAATTCACAACCTCGACTACCATTGTTAGACAGGCTATCGTCCGTCTCTTTATCTAAGAGACCGGAGCGCCCACAACAAAGCCTACCATCACTAAGGCATCTGCAATTATTACCC tpg|BK006944.2|:93797-95011 7X148= 219S3=7X 
 tpg|BK006944.2| 642804 + tpg|BK006944.2| 643287 - INS TTTAACGTTGCCTCTGTTCTTTTCCTATTAATTCTATTAGATAAGTTTATTTCCATCTCATATAAAGAAGAACCTGTCGAGGTTATATGATCTCTTTTCCGTCTTTTTACCGATTCTGGTTAGTGTATGCTTCATTTGAGTTTCTTGCACTGCTTTGCCGACCAAATATGGAAATCATCTATTTTAACTCTATTATTGAAGAGGCTTTTCCTGGCACATAT tpg|BK006944.2|:642348-643743 7X182=18S 1=204S 
 tpg|BK006944.2| 507812 + tpg|BK006944.2| 508226 - INS CGAAAGAGGTTAATGTTGACGACGAAAAGGAAGACAAACTTGCACAAAGACTAAGAGCATTGAGGGGCTGAAAAAACATGCTAACAGGTCATGCATTTTTAGTTCATCATTACGTTTCCAGCTATGTTATGTATGTATGACCACATATGCTGTACATAAATTGTATAC tpg|BK006944.2|:507462-508576 7X94=32S 3S1=235S 
 tpg|BK006944.2| 614608 + tpg|BK006944.2| 614694 - INS TTTGTGTCAAGACAGAGAAGTGGGCTGCTTCTCCCCTTTCAACACTCCCCTCCCATGGCTGAATACTCAGACGTTTTCTGTGGTGGAAATGGCATCAAAAGTGCCACTGGCTGGCGAATCCAGACTATTTTGTGTCAAAGAAACATGCGTACCTGCACAATAAAAAGA tpg|BK006944.2|:614258-615044 7X9=75S 79S5=7X 
 tpg|BK006949.2| 464140 + tpg|BK006949.2| 463917 - INS CAGGGTTTGGTCCCAAGAGTGAGATTAGTGTAGTCCTGGACGTTAAGGTTGTTACGCCAGATGCCGCCGCTGAACAGTTCGCAAGGGACTTTCCCTTGAAGAAGGTTCCGGCTTTCGTGGGTCCAAAGGGTTACAAGCTAACCGAGGCAATGGCGATTAACTATTATTTAGTAAAGCTTTCACAGGACGACAAGATGAAGACTCAACTTTTAGGTGCCGACGATGACTTAAATGC tpg|BK006949.2|:463433-464624 42S82= 67=58S 
 tpg|BK006944.2| 417222 + tpg|BK006944.2| 416596 - INS CAGTACTCAGACCGCTCCCAATAGTCACAGTACTAGTATCAGATGACAAAACTCGTAAGGTTTTAGTCAGTAATGAGGTAGTTTTCGAGAATTTCCCATGGTTATTTACTTGAGCATAATATGACCAAGTCTGTACCAATTGAGCACCAAATCCTCTTTGGAAGAACACTATTAGAGGTTGGTAATCTTTGGAGAGAGTTTCATCTTCGACTGCACTGATTATACTTTCTAGTGTTTCTAATGTACCG tpg|BK006944.2|:416086-417732 8X11= 13=1X219=7X 
 tpg|BK006944.2| 206163 + tpg|BK006944.2| 206703 - INS GATATAGATTACTCTACAATTTCTTTGTATACAGCGGGAAATTGACACTTCAAAGTTCCTCTCATATCAACAAACATTAATACAGTTCCTGAAAATGTATTCTTGGAAGTCAAAGTTTAAGTTTGGAAAATCTAAAGAAGAAAAAGAAGCCAAACATAGTGGGTTTTTTCA tpg|BK006944.2|:205807-207059 7X6=79S 81S5=7X 
 tpg|BK006949.2| 522269 + tpg|BK006949.2| 522864 - INS AGACAATGGTTACGATATCAATTACATCTCTAAAATAGGAGACAAAATAGATTCCAACAAGCCAATTTTTCTCTTCGCGCCAGAGTTAGGTGCAATTAATTTACATGCTTTATCAATGTCCCTCCAATCGAAGAATCTTGGAGAAATAAACACCGCCTTGAACACCTTGTTGGTCACAAGCGCTGACTCGAACTTAAAAATATCTCTGGTCAAATACCCTGAATTATTAGACTCCTTGGCAATACTCGGCATGAATTTACTGTCAAATTTGTCACAAAATGTTGTTCCATACCATCGAAACACTTCTGACTATTATTATGAGGATGCTGGATCAAATCAATACTATGTTACCCAACACGATAAAATGGTTGATAAAATTTTTGAAAAGGTAAACAACAACGCTACACTTACACCGAATGATTCTAACGATGAAAAAGTCACTATCCTGGTAGATTCTTTAACAGGTAATCAATTGCCCACCCCTACTC tpg|BK006949.2|:521279-523854 7X183= 244=7X 
 tpg|BK006944.2| 118867 + tpg|BK006944.2| 119148 - INS GGTTCACATTCGCATTCGCACTCACACTCACATGCGGATTCGCATTCGAATTTTAGCAACGATCATGATTTAGAAAATGCTCCCTCTGAGCATGGTTATGCAACATCTTCTTCCAGTGTTTCTGAAAATGACCCGTTGATTACAAAGGATAGCGATAGACCCCAAATGAAAAAGAAAATGTCCCTAATTGACTTATTAACCAGAAGGAAATCAGAAGGCGAGTGT tpg|BK006944.2|:118403-119612 7X5=140S 113=7X 
 tpg|BK006944.2| 222933 + tpg|BK006944.2| 223141 - INS CAAACTTGTCTAACTGTTCCTTACGCGATTTAGCACCTAATTTCTGCAGCGTATCATTTTTTTCTTTATACTCCTTGTCTTCTAACAATTCGCTCTCACTCTTTGATTCCAACCACTCCATAAGTTTGATTTCATTACCATAGCCTTCATCATTTTCGTATGGAGTTTCCAAGACAATAGGGATACCCTGCAGGTATTCAGAGTGCGCGATCATTCTAAACACATCTATAC tpg|BK006944.2|:222457-223617 7X150=23S 6S1=48S 
 tpg|BK006944.2| 220007 + tpg|BK006944.2| 219780 - INS TGTTATTTGTGACCTCATTTACTCAGAAGAATTTCGTAAATCGGTTGTTATAGAACTGTTTTATTGTTTAAAAGAGCTTGTTATAGTAATCTAAGTGGAAATACACTAACAGTAAATAGGGCGTGTGGCGTAGTCGGTAGCGCGCTCCCTTAGCATGGGAG tpg|BK006944.2|:219444-220343 7X4=166S 81=7X 
 tpg|BK006949.2| 812789 + tpg|BK006949.2| 813286 - INS GGGCATATATATCCGAGAGTACTTGTGGCTCGTTGATCTTGCATTTAACATTAATGCCCTTGTTCAGAAATCTAGATAAATACTCCATATTGGAGATGGGCAATGTGGTGATGGCAGTTTTATTAGTTTTGATTTGGATGGTCTGCAATTCAAATTTTTTAGTTTTGGCCATTGCGGGGTTCATTGTGGTTATTGAAGGGTCTATGAATTCTTTAAGTTTTTTCCCGGTTATACTAAACGGTAAGACGCTTTTACCATTACATGAGGTACCCTCAGCAAACATAAAATTCACGGTATTGCCCAATTGAGAT tpg|BK006949.2|:812153-813922 7X189= 292=7X 
 tpg|BK006944.2| 660165 + tpg|BK006944.2| 660611 - INS AACCTGATGACACTATTATCTTTTGCATATTTTGTCGACTCGTATCATGTACGCGCTGCATATGAGGTGCGGCGCTATCTGTTAAATATGTACTAATTTGAACCTGCTGCAAAGGAAATGTGGCACTACTTTTACTCGCATGTTAACTTTCACCTACTATATATAGAAAAAAGGGTGTTGCTTTCAATCGCCGACTAATTTGCTCAAATACTCTTTACACAAAGGAAATTGTGTATCAGTAACCCTTACGGTTTGTTTATGAAGGAACTTTGCTCGTCCTACACCACCGGATCTAGGTACTCAATTTTTTGATGATTTTGCACTTGTGCTCATATCCTGTCGACAGGCACCGCAT tpg|BK006944.2|:659441-661335 11S96=1X76= 178=7X 
 tpg|BK006944.2| 208111 + tpg|BK006944.2| 208523 - INS AGCTCATGATATGCTTAAATATTTCTTAAGGATGATTCCCTCCTCGATGGGATTCATAGATACATATTTGGCCAAATTTTTCCCAAATAAAAATGATACTCGGAGAAAGTTGGTTAATTACACTTCAAATTTGCTGAAATTGAGAGGCTACTGCTCTGAGCTAGGA tpg|BK006944.2|:207765-208869 7X1=2I108=34S 4S1=129S 
 tpg|BK006944.2| 256469 + tpg|BK006944.2| 256701 - INS GAACTACTCTTCCATTGAACAGCAACACCTGCAAAATCGGAGCTGCAAAATTATTGATTGGATGTGGCAAAAATAGGAATGGGCGATCATAATCTGCCGGATTTTCAGACATGTTTGAAGTTTTCTGTTACAGCTAAAAAGAGCTTTCTATGTATGTATAG tpg|BK006944.2|:256133-257037 7X6=145S 141=7X 
 tpg|BK006944.2| 265208 + tpg|BK006944.2| 265272 - INS AAGAACAGGTGTGTGTGCTAAGTAAGAAGAATTATTACATTTACCCAACATGAGGATGGAAAAAACAACAGACAAACCACTTTCTGCAGGAGATATGAACGATGAATATTCTCGGGGTCCAATCG tpg|BK006944.2|:264944-265536 7X5=57S 59S4=7X 
 tpg|BK006949.2| 871674 + tpg|BK006949.2| 871797 - INS GCTTGTCAGGAGAGACTGAATTCCACTCATTCCAATTGAAGGCTCTCAAGGGAATCAAGTCATTTTTTCCAGCTCCTTTATTGTTATTAAAATTACAAGAACTACACCCACATACATTTAAAAAATTCCAATATTGTACCATAATATCCTCCTCGACAGGAAATATTTGTTTTTGCGTCACCGAACGATCGACAATAGT tpg|BK006949.2|:871262-872209 122S119= 100=7X 
 tpg|BK006944.2| 224160 + tpg|BK006944.2| 224005 - INS TTCAAAGTCTCCATATTTACAATGATTTCCAACATGTAAAGAAATGAAGAAAAAGAAACCAGGTAAGAATGAAAAATTCCACGTTCAAGTTCCCAGAAAAACTGGCAAAAAAAGAGAAGTATTAGATGAAAAAAGTTCGTGTATACAAATATCTATGTTACATATATGCCAAGGTGAAGGACCAAAAGAAGAAAGTGGAAAAAGAACCCCCTCATCTTCTTCCC tpg|BK006944.2|:223543-224622 19S95=5S 107S5=7X 
 tpg|BK006949.2| 604360 + tpg|BK006949.2| 604378 - INS GCATCATCCCGCATGTCATTCATCTCCAAGGTGCTCCTGCATATATGTAATAATCATGATGAAGAATACGTAGGACAATTTGAGAGATATGAATAACGGGAATTTTACAATTTGACGGATTATCGGAGGAAAGCAAGTCCAAATCATCATCACATAGTCCATCTCCATTATCCTCGTCAATTTTTCTGTTCGTTAGTGTCTCCTCAGATGGAGTACTTATCCTACATGCTTTCGGATCAGTGCAGCTTTTCTGAACTTCGTGAAGCCAATAGTTC tpg|BK006949.2|:603796-604942 7X185= 5S253=7X 
 tpg|BK006944.2| 451542 + tpg|BK006944.2| 451427 - INS GAGGGCAGGTGATGACAACCTCAGTGGGCACTCAGTGCCTTCAAGCGGATCCGCACAGGCAACTACTCACCAAACTGCACCAAGGACTAATACGTTTACTCTGCTTACATCACCGGATTCAGCGAAAATATCAAAGGAACAGTTAAAGAAGTTGCACTCTAATATAC tpg|BK006944.2|:451079-451890 7X3=1X127=15S 11S1=202S 
 tpg|BK006944.2| 645161 + tpg|BK006944.2| 645415 - INS GCATTGAGACCCTATATTCCCCTCATCTATTCCAAATAAGAATCATATAAAGAATTCACTAGGCACAGATAACTGCTGATTTATAGACATAATCCCTTCGCATCCACGTTAGCATGATTGGTGACACGCTTTCTGAGCATTAGCTTGCGATAGGTTTCCAGCAT tpg|BK006944.2|:644819-645757 7X6=76S 78S4=7X 
 tpg|BK006944.2| 270936 + tpg|BK006944.2| 270355 - INS CTCCCATCCTTCGGCTTCCTTGTTGTTTTCATAATCCTCGATAATAGTGTTGGCACCGTATTCTTCCCTCCATCGTTCAGTTTCTACAAACATCTCAACGCTAGCATTGATATCAAATTTCCTTGCCCGTAGAAATCGCAATAGCGTAGAA tpg|BK006944.2|:270039-271252 7X4=215S 133=7X 
 tpg|BK006949.2| 273231 + tpg|BK006949.2| 273439 - INS TTTTCCTGGTGATGAGAACTTGGCTCTCTTTGTTTGTAGCCAAGCTGGATGGACAAATAGTCAAAAATATAATTGCTGGTAGAGGAAGAAGCTTTCTGTGGGACTTAGGGTGTTGGTTTTTAATTGCTGTCCCTGCTTCTTATACTAATAGTGCTATTAAGCTACTTCAAAGGAAGTTGAGTTTAAACTTTAGGGTAAATTTGACACGTTACATCCATGACATGTATTTGGATAAAAGACTAACATTTTACAAATTAATTTTTGATGCAAAGGCGTCCAATTCGGTAATCAAGAATATCGACAACTCCATTACTA tpg|BK006949.2|:272587-274083 7X186=50S 2S1=156S 
 tpg|BK006944.2| 243629 + tpg|BK006944.2| 243617 - INS GTCTCTGAAGACACCACAGCAGCAGCAAATTGGTAACCTCTACCCAATAACAATAGAGATTTTTGATCCTTTAATTCAGTCGCACAGAGCTTTTTTATTCTTGGTTCCAGCTTTAATACCTGCTTAATTTGGCCCGGGATTAACTTCAAGCCTTGAATGATTTCAATTCTTC tpg|BK006944.2|:243259-243987 7X296=4S 151=7X 
 tpg|BK006949.2| 668187 + tpg|BK006949.2| 668164 - INS GGGTTTCATATTCAATATTACAACTTGAGTTACAAGAACATTTACTTTTCAACAATCTGATTGAAGAAATTCACGACATTATGTACTCCAAATCTAACAAAACAAATTTTACTCGAGTAACCAATAATGATATATTCAAAATCATAAGCATTTCACATAATGGATTTACGAGTTTAGAAAATTACCTGTACAACATAGTCAATATTGATATTATGGAACACTCAAAAACGATAAACAAGAACC tpg|BK006949.2|:667664-668687 25S169= 4S224=7X 
 tpg|BK006944.2| 337426 + tpg|BK006944.2| 337496 - INS ATTACCACTGTTGCTGTGGTTGTTGTTGTTGCTGTGGTTGCTGTGGTTGCTGTGGTTGCTGTGGTTGCTGTGGTTGCTGTGGTTGTTGGGATTGTTGTTGTGGTTGAGGTACAGTATTAGCTTGATCTTCTGGAGGCTCTGAAATAACAGCACTAATTTCAACCTTTTCTTCAACAACTGTAACTTCTTCTTCTGGAGCAGCAACATTATCTTGTTCTTGTTCCAGCTCTTCCGCTGTCTGTTCCTCTTCTTTTACTTGTTCCTTTTTTTCAGCTTCTTCTTGGAC tpg|BK006944.2|:336840-338082 7X5=17S 269=7X 
 tpg|BK006944.2| 281942 + tpg|BK006944.2| 281979 - INS TTGAATAGGATCGTTTACTTCTACGTTCAGGTCGGAGTCTCCTTCCACTTTTGATGTTGCTTCCTTTTGCTTTTGCATTTTCATGTGCTTGAATTTTTCACCAGGTAGGACCACCGGCTTTGCGTCTTTCTCCTTCTTCTTCATTACTTCTAATGTACTAGATGTTTCATCATCACGTTGCTCCGGGTCTAATT tpg|BK006944.2|:281540-282381 7X178= 97=7X 
 tpg|BK006944.2| 664450 + tpg|BK006944.2| 664904 - INS ACGAGACCGTAGGGACATATAGCACCTTAGAAATAACCTTGTATGAAATCTTTCATTATTTCCTGTTTAGACACTTGCGTCAAGGTATTTTTTTTATCGTGGTGTTGAATGTGGTAACCCAATAGCATAATATGAGTAATGCTTTAGTATTGTTTCAGAGCTGTTTTAGATAAAGAAAACACATAGTAGCAAACCTCTAATCCGGTAGTACTTAAGAAACTATAGTTTCTATGTAC tpg|BK006944.2|:663964-665390 7X63=55S 6S1=264S 
 tpg|BK006949.2| 896268 + tpg|BK006949.2| 896350 - INS GTGTAAGTCACTAGTATCTTGCCGTTAACCCTGTCCTTATTGCAATATGGTCTCAACCAAAAGGGCAAGGCCATAAGCTTTGAACAAATGAAAAGAGATGCGGCCGTATGGTGTGAAAATCTGGGTGTACCAGCAACAGTGGTAAAGGACGATTACATACAACAGTTTATCAAACAGAAA tpg|BK006949.2|:895894-896724 12S42=43S 83S7=7X 
 tpg|BK006944.2| 443199 + tpg|BK006944.2| 442718 - INS GTTTCCACCGCCAAAGCGTCTTCAGATTGTCC tpg|BK006944.2|:442640-443277 7X10=6S 12S4=7X 
 tpg|BK006944.2| 27290 + tpg|BK006944.2| 27729 - INS CCAGATCATATTCAACCATTTTTGCAAGCATTTTTTTTATGGATTCAGATGCATTTGTCTGAATTGCAGCCATGTATTTCAATATTGTAGCCAGATCATATTCCTTAGTTAATGACCCAATTAACTGTATCCCTTTTGTGTTAGCTGCGACTTGCGCTTTTAAATCGCTTATGTTATCACTAAATCTTCTTGAACCTGAGCAGCCTGGGTATTTGCCTGGATCTTCTA tpg|BK006944.2|:26820-28199 7X156= 214=7X 
 tpg|BK006944.2| 481098 + tpg|BK006944.2| 481456 - INS AGATGCTAGGCAGTAGTGACGAAGATGCCTTTCCCAAAAGCCAATCATTAAATTTCAATAAGAAACGACCAATACTTAAAATTAATGATAACGTCATACAATCAAACAGCAATAGTAATAACAGAGTTGATAATCCAGAAGATACAGTGGATTCTTCAGTCGATATTACAGC tpg|BK006944.2|:480740-481814 7X66=1X89=5S 7S1=30S 
 tpg|BK006944.2| 169170 + tpg|BK006944.2| 169210 - INS GCTGTAGTGGTTTGTGTGGCAACCCAGGCTGTAAAGTGTCAGCAACCGTATGGGCAACAGCACGACCAAAGACAACAAGATCCAACAAGGAATTGGCACCTAATCTATTG tpg|BK006944.2|:168936-169444 7X5=50S 51S4=7X 
 tpg|BK006944.2| 183066 + tpg|BK006944.2| 183714 - INS CCTAAGGATACGAGAGGCTGAATTCCTG tpg|BK006944.2|:182996-183784 7X10=4S 14=7X 
 tpg|BK006944.2| 447388 + tpg|BK006944.2| 447292 - INS AAAAGATATGGAAGAACCAGTGT tpg|BK006944.2|:447232-447448 7X4=7S 12=5X2S 
 tpg|BK006944.2| 28528 + tpg|BK006944.2| 28547 - INS CATTTGTCTGAATTGCAGCCATGTATTTCAATATTGTAGCCAGATCATATTCCTTAGTTAATGACCCAATTAACTGTATCCCTTTTGTGTTAGCTGCGACTTGCGCTTTTAAATCGCTTATGTTATCACTAAATCTTCTTGAACCTGAGCAGCCTGGGTATTTGCCTGGATCTTCTACGAAA tpg|BK006944.2|:28150-28925 7X7=84S 87S4=7X 
 tpg|BK006944.2| 458780 + tpg|BK006944.2| 458508 - INS CTTTGTATTTATTTCATTGTCATCCACATCCAGCATTGGTTTTCCATTAGAATTTCCAGCTGGTCCATGACTTGTTTTGAAATTAATTTTTTTAACTTGCACGTTCCTCGAATCAGAATCATCATCCGAATCATCTGAGGAAGAGCTATCCAATGAAGATTCAAGTGACATGGAA tpg|BK006944.2|:458144-459144 7X87= 189S3=7X 
 tpg|BK006944.2| 365697 + tpg|BK006944.2| 365351 - INS CCTCAAAAAATAAAAAAAGTCAAAATAAGAACACATCAGTTAGGAACCGTGCTTGGAGTTTTGAGACTGGAGTATTGTCCATCCAACATATTCTGCTCTTTCACCATAGACTTCGTTGGAAATCGCCTCTCCCTTGTACTATATTGTGCAGAAC tpg|BK006944.2|:365029-366019 7X5=68S 77=7X 
 tpg|BK006944.2| 291225 + tpg|BK006944.2| 290783 - INS CACGATAGTATACGGTTTATGGA tpg|BK006944.2|:290723-291285 7X4=7S 7S5=7X 
 tpg|BK006948.2| 159673 + tpg|BK006948.2| 159381 - INS GATAGAGCCCAACTGAAGGCTAGGCTGTGGATCCGTGTGGAAGAACGATTACAACAGGTGTTGTCCTCTGAGGACATAAAATACACACCGAGATTCATCAACTCATTGCTGGAGTTAGCATATCTACAATTGGGTGAAATGGGGAGCGATTTGCAGGCATTTGCTCGGCATGCCGGTAGAGGTGTGGTCAATAAGAGCGACCTCATGCTATACCTGAGAAAGCAACCTGACCTACAGGAAAGAGTTACTCAAGAATAAGAATTTTCGTTTTAAAACCTAAGAGTCACTTTAAAATTTGTATACACTTATTTTTTTTATAACTTATTTAATAATAAAAATCATAAATCATAAGAAATTCGCTTATTTAGAAGTGTCAACAACGTATCTACCAACGATTTGACCCTTTTCCATCTTTTCGTAAATTTCTGGCAAGGTAGACAAGCCGACAACCTTGATTGGAGACTTGACCAAACCTCTGGCGAAGAATTGTTAATTAAGAGCTTATTTACCGCTTTTACGTAACGCCCTACGCTTGTTCCATAAGCTTTGTAAATCGTCTACAGGAGTGCTCTCGTGTAGCTGTATTGTATCTTCAATTGGATAGTCCGTAGTGATGCTTTTCGGAGAATCGCTATTAACTCCAGCAAGTTCGGCCATTTTTTTGCCGTTTTTTGCCTTCTTCGCTCTATGGGGCAGAGACATCTGTCTTAGGTTCTCGTGTTCTTGTTTGATTCTTTCATGTAGGGCCTGCCTGGCCTTTGCCAGGCTCAGTGAGTCTACTTGACCCTTAATAAAATCCCTGTGCACCTTGACTGTTCTTAAGTGTTCACATAAGGACAATTTTTTCGTATATCCAAGCGGATCATATTTACACGGAACTTCGATGTATCCTTTTTTCTCTTCCAGAAATACGAATATTCTGCTCAGATCATCCGG tpg|BK006948.2|:157495-161559 7X486=216S 673S4=7X 
 tpg|BK006944.2| 255782 + tpg|BK006944.2| 255462 - INS CTATAAAA tpg|BK006944.2|:255432-255812 7X4= 4=7X 
 tpg|BK006949.2| 382565 + tpg|BK006949.2| 382713 - INS GATATATAAATCATGGGCCCACTGATATATAGAAGGCTAAATAACGAGAATCATATATACTGTAACATGACACCTGCTGATTTTTACTGATCGTAGCCATTCGGCTCATATTACTTCATGTCCCTTTTTTAAATCCCTCGTTCCCGGAGAGTGGCATAGCATGTCCGATAGCGTACGCCAACCTACAGAATCAGGGGATCAGATTTCCTGAAAGCAACTTATCCATCAGTTTCTTTTTATAATGCCATAATGACAGGTG tpg|BK006949.2|:382033-383245 7X8=8S 237=13S 
 tpg|BK006949.2| 94720 + tpg|BK006949.2| 94728 - INS GATGGTAAAACTTTCTACTTTTTTTGACAAAATTGTCGCAGAACTGTTGCTAGCTGACGTCTTAGTCTTTAAATGACTTGGCGACGCTATGTTTAACGAAGAGTTGATTTTGGAACTTGACTGCGGTCTCAGAGGTGGAGTCACATTGGTGCCTAGGTTTTCAACATAACGATTTAGATAAGAATTATTATTGCCTGGTTTCGAAGGAGAGCCTGAATATGCTGTCATTGTT tpg|BK006949.2|:94242-95206 185S80= 218=7X 
 tpg|BK006949.2| 879618 + tpg|BK006949.2| 880170 - INS TTAGATCCGAGTTTCCGCGCTTCCACCATTTAGTATGATTCATATTTTATATAATATATAGGATAAGTAACATCCCGTGAATCAAGCTGATAAACAGTTTTGACAACTGGTTACTTCCCTAAGACTGTTTATATTAGGATTGTCAAGACACTCCGGTATTACTCGAGCCCGTAATACAACAGTGAGCTATTAAAAGAGCTTAAGTATTACAGAGTAATATCAATCATCAATCTTGGATCTAAAGTAATCGTCGAGACATTTATACACTTAAGTGATTCCTCTTTACAAGCGGAGCTTACTC tpg|BK006949.2|:879002-880786 7X241=22S 4S1=68S 
 tpg|BK006949.2| 428959 + tpg|BK006949.2| 429720 - INS CCATCTTTGATCTTACAGATGATATGCTGTTCCAGGCCGGTGTTGACGTCGATGAGAAGGGCCAAGGCAAAAACGAGGAAACATCAGGAGAAGGAGGAGAGGACAAGAATGAACCTTCTTCCAAAAGTGAAAAATCTAGAAGAAAAAGACAAACTTCTACAGATATTAAA tpg|BK006949.2|:428605-430074 7X8=77S 79S6=7X 
 tpg|BK006949.2| 885954 + tpg|BK006949.2| 885877 - INS GCGCCACAACGTAAAATTTCTTTGCCAGAGGCATTGCGAAAAGTCGAATTGATGAAAAAATCTAAAACCGAGCCTGTTTTAGAGTCCTCAAACGAACTGAGCATAAACGCAAAATTAGACGCAATAATTGCCTCTAGAAACTTAAGAGCATCTAATACTCTACCAGAACTTAGCGGTGTTAACACTAATAT tpg|BK006949.2|:885481-886350 7X4=91S 84S5=1X6=7X 
 tpg|BK006949.2| 884641 + tpg|BK006949.2| 884345 - INS AAGACCAGGAAGAGCCGATATACCCTCCTCCTCCTCTTCTTCATCACCACCGCCTTTGCCCACAAGGCGTGATCATATCAAAATCACAGATGGGAATGAAGAGAAACCGCTTCTTCCAACAAGGCCTAACAAAGCAGAAGTTACAGAAAGTCCGTCATCAAGGTCAATAAAACCGGATGCTGTGGTACCTGAGCGCGTTAAGCCTGCTCCACCTGTCTCACGCTCTACAAAAC tpg|BK006949.2|:883865-885121 7X5=336S 117=7X 
 tpg|BK006949.2| 937430 + tpg|BK006949.2| 937430 - INS TTCTAGTATTATGAAGAATTCCAAGTTAATCGACGAAAAGCGTTTGGAAAGGAATTATATAAACGTAAACATGAAAAATATTCATCGAATACTCCACATCGATCGTATTACAGTGTTTTAGTAAATGTTTGTATTTGAATCAAAGTTTCAGCATTTGTTCTACACTGATAAAATCATGGTTCTAGTATAGTGAAACATACGCCCAAGTTATCCTAGTACAAGACCGCCATATTGTGCTCATAATCGGGAACAATGAAAATAACACCCTAACAATTGCTGAAACTTGTCGTACGCGATCCCTAATTACATTATCAAGCATTCAGCATTGGTCAATACCTCAATACCTCGACAAGAAAAAAGAAATAGACACGTGTATGTCAAGGCATTAAGAAGGGTATCAGGCCTAGTGCTCGCCTCTTGCCTTCCCAATTTGTTGAACATCTTTGACATATAATTTGATTTTGAAATAGTTATTGGACTTCCATTTTAAATAAAGGCTCTATCATTAACTATACAGAATATACTAGTAACGTGAATACTAGTCGATAGACGATAAATTAATACTTTTTCCAATAAAATCTAAACGCATGCAAGTACATAAATAGGCGAAGGTATCTGACCGTAATAATCTTCACGCCATCTATATAAATAAATGAAAAATTCGGCTTTTAACTTATATATTAACAATAAGAAAGACAATGTTGCGCTGTGCTTACA tpg|BK006949.2|:935982-938878 7X6=148S 695=7X 
 tpg|BK006949.2| 329861 + tpg|BK006949.2| 329880 - INS CTTAATAACCTATACTATTCTGTGACTGTTATTTATTTACCCTCGTAATATTAAAAATGTCCTATACAATTTCTGTAATAAAACCTAATTTTTTTAGGACCCTTGAGTGTTACCCTGCTCATGTTTTTATTTTTGTTTTAGAGAAATGTAAACAACAGTTTGGGAA tpg|BK006949.2|:329515-330226 7X5=78S 78S5=7X 
 tpg|BK006949.2| 396318 + tpg|BK006949.2| 396908 - INS AGTAGAGACTGTGCAGTTTTTTTTTGAAAACTTGCTTTCATAGACGACTCACTTTTTTCAGTTTGAGATTTCGCGCTCCTCTTATGAATATATTCCTTTCGTGGGATATCTTCAACGT tpg|BK006949.2|:396068-397158 7X3=164S 59=7X 
 tpg|BK006949.2| 711927 + tpg|BK006949.2| 711961 - INS AGTTTAGATATTTGATAATGGACCCATTTTCATTATTGTTTGCATCTGTTTCTTGAAATCTAGCAAGGTGAACTTACCCTTTTGGATGTTTTCCATTGTGGCTTTTGCATCTTCCTTGTTGGAAACGGTTTGTAATTGCTCAAAGAGACTCTCTATATCACCAATACCCAACAGTTTAGATATGAATGACTTAGGCGAGAACTTTTCCAAATCATGAATGTGCTCACCTGTACCAATAAAGATAATCGGAGTGTTTGTGGCTGCAACGGCCGAAATTGCCCCACCCCCTCTAGCGTGGCCGTCCATCTTGGTTAATATAATGGCACCAAAATCGGACGATTCTTTGAAAGCCTTGGATTGTTGCTCTGCAGCTTGACCAATGGAAGCATCTAAAACCATGATAGTTTGATTAGGCTTGATGACATTGGATATTTCAATC tpg|BK006949.2|:711035-712853 7X195= 220=7X 
 tpg|BK006949.2| 619050 + tpg|BK006949.2| 619112 - INS CTTTGGAGTGTATGATGAAAATATCATGCATGCTTATATAAAAGCTTTTTTTTTTCTATAGGGTGACATTTAGGAGCAATAATTTTTACTACAAGCTTTTTTTGCACCTTATATAGTAGTGACCTTGAAATTGGTCTTTTGCACCAGCGTACTTTAATTCCACTAAGTACTGTTTAGCAGCCTGTTTTCCAGAGCCCACAAC tpg|BK006949.2|:618632-619530 7X15=19S 3S187=7X 
 tpg|BK006949.2| 470636 + tpg|BK006949.2| 470707 - INS AAACCTGTTATCGATAAGTCTACGGGGTTGGCTAAAGGTACGGCCTTTGTAGCCTTCAAAAACCAATATACATATAACGAGTGTATCAAAAATGCGCCTGCGGCTGGCTCTACCTCTTTATTGATAGGTGATGATGTCATGCCTGAGTATGTGTATGAAGGTCGTGTTCTGTCCATTACTCCAACGTTAGTAAGAGAGGATGCTGGAAGAATGGCAGAAAAGAACGCCGCCAAAAGAAAGGAGGCCCTAGGTAAAGCGCCAGGCGAAAAAGATAGACGTAACTTATATTTGCTGAATGAAGGTAGAGTTGTTGAAGGCTCAAAAATGGCTGATTTGTTAACCAACACTGACATGGAGATCAGAGAAAAATCTTACAAATTAAGAGTGGAGCAACTGAAAAAGAACCCATCTTTGCATTTGTCGATGACTAGGTTGGCTATCAGAAATCTTCCTAGAGC tpg|BK006949.2|:469706-471637 7X152=1X6= 229=7X 
 tpg|BK006949.2| 568649 + tpg|BK006949.2| 568090 - INS CCTTTGATCTCTTATTATACCCCTAATGAATTCGTGGTCTCTCGGATCACTGCTTGAACTCAACAGCTTACCATTACAGGAATCTGTTCTTGCAATAACCAAATTTTCTGTCCCCATGATATCCCATTGAAACCTGGTGGAAATCAATCTCATAAGATGTGTTGCTGTGGGCACCAAAACAGCCCCACTTAGATGGCCACACCTTTTGCCTCCCACCATCTGATCTTCAAGATGAATACCAGCAGCCCCTTTCTCCGCAAACAACTTAGCAACTTTCATTACAGTCGTTGGGCCACCGTGACCCATGTCTGCGTCCGCGATAATTGGTTTTAAATAATCAACAGGAGTAGAAC tpg|BK006949.2|:567370-569369 7X5=148S 177=7X 
 tpg|BK006949.2| 269344 + tpg|BK006949.2| 269981 - INS CGACTGCGTCGAGCACCTCTGAAAGAAGTTCAAGAACAGATGCCTTTTACGATATCACTACAGCTACACCAGTTGTGACCACTGATAATAGGCGCAATAAAAACAATAATCTGAAAGAGTCTGTTTTGCCCAGATTTGGGACTCAAAGGCCATGGACTGGCAAAAGGACGTATACCACGTCCCGCCATGGCAAGAATGCTAGGCGTTCGTCTAAAAGAGGTCTGTTCAAAAT tpg|BK006949.2|:268866-270459 7X41=1X138=23S 2S1=154S 
 tpg|BK006949.2| 321566 + tpg|BK006949.2| 321715 - INS TTTTACAAGTCACTTTCATATAGAAAGTTGGTATATAAAGTGTCAACTAAGAGAGAAATAGTTCGAACCAGGTGTATTTTAAATCAACTATCGGGAAGTATGGACTGGTGGTATAATCGAATTACATAGTCCTTTTACCTTCATTAGTAGTACTTAAGTGTCACCCGCCTGGGGATTTTGCTCTCATAGAAGTAAAAGGGTAGTGCTATGGGAGCACATTAGGT tpg|BK006949.2|:321104-322177 7X128= 210=7X 
 tpg|BK006949.2| 860252 + tpg|BK006949.2| 860285 - INS GCTATATCCGTGACATGCGATCCAAGTGACTATCCAACATATGATTATATTCAATCGCACTTAAATGCATTCCAGAATGCAAACTTAACTACTTGGGAAGATGCTGGTTACACGTTCCCTAAGAATATCCTAACTGGTAAATGTACTAGCTCGAAGTTCAAGTTATCCTCTTAAGCGGGTATTTTGATGGTAAATCTCCAA tpg|BK006949.2|:859836-860701 7X3=97S 96S5=7X 
 tpg|BK006949.2| 829733 + tpg|BK006949.2| 829776 - INS AACTACTGTATGTTTGCTTGTGCATATGGTATATTCACCGATTCATTGTACGGTGTCTTTGCCAACTTCATTGAACCATTGGCATGGCCACTAGTTTTGTTCACACTGGACTTTTTGAACTTTGTGTTCACTTTCACTGCCGGTACAGTGTTGGCCGTTGGTATCAGAGCTCACTCATGTAACAACAGC tpg|BK006949.2|:829341-830168 7X137=28S 1S1=13S 
 tpg|BK006949.2| 157507 + tpg|BK006949.2| 157547 - INS ATATAGACAATCCCAGCATCAAGATTCCTCCCGAGATTGTCATTTCAAGGAATCTGCCCATGAAGTTTTTTGGGCTAAGTGAATCCACTAAGAATATCAACGGATGGCTGAAGTTGTTCTTCGCAAAAATAAAATTTGATAGGGATAATGATACTATCGTGGAC tpg|BK006949.2|:157165-157889 7X5=77S 77S5=7X 
 tpg|BK006949.2| 401064 + tpg|BK006949.2| 400932 - INS GTGTAAGTTTTGCGGATTCTTTGGCTGAATTGATTGCCATCAACACGCGATGCTTAGAATCTTCTAATGGCTTCTTGGCCAATAGTTTGTAAGAGTTGTTCATGGATTTGAACATTTTATCATAGTATTCGCCGTACACTTTTTCTGCTGTTTCAACACCAAACGCATGTGGACCGGCTTCTGTTTCGCCTTGAACCACAATTGCTACGTTGGGTAGTTTGTACTGAGGTAACATACCTACATCCACAAAGGTAGCCAGTAGGCTTTGACATTGAGTCCTCAGAGCTTTTAAGCTAGGTACTAGC tpg|BK006949.2|:400308-401688 7X203= 153=7X 
 tpg|BK006949.2| 286165 + tpg|BK006949.2| 286144 - INS TTTTGCTGTTCTACACTCATTCTTTCGATTGTTTTCAATTGCTTTTTTAGGAAGTGCGGCTTTGTTTACATAAAAGGTGTGCGGCATTTTAATGCAATATGAAATTTAAAAGTATATGTAACGATAGCACTATTATTTAGGGTTCCTGAAATGATATACTTTATGGATAGACATTATCTGTTCATTGAGTATACAGT tpg|BK006949.2|:285736-286573 7X140=32S 2S1=173S 
 tpg|BK006949.2| 751765 + tpg|BK006949.2| 752032 - INS TCTATCTTAGAAGATAGACAATGATATCTTGTGATAGTACAAGATGAGTTCGAATTCAACACCAGAAAAGGTTACTGCAGAACACGTTCTGTGGTATATTCCCAATAAGATCGGTTATGTTCGTGTTATCACCGCCGCCCTTTCTTTTTTCGTTATGAAGAATCATCCTACGGCCTTTACATGGTTGTATAGTACATCATGTCTACTGGATGCGCTAGACGGAAC tpg|BK006949.2|:751301-752496 75S150= 8S196=7X 
 tpg|BK006949.2| 748809 + tpg|BK006949.2| 748276 - INS TTAGGCCTATATTGAAGCATGAAAATACGCTTAGAAGAAGTAAAGAATTTGGAATTTCCTGCTTTCACAGAAAGGTCTAGCGAGGATAGAAGGAAAATATATCATAACATGAGGAAGACAGAAATTAATTACGCTAACTCTATGGTCGGTTCGCCTGATTATATGGCCCTAGAAGTTCTGGAAGGTAAAAAATACGATTTTACAGTGGATTATTGGTCATTAGGCTGTATGCTTTTTGAAAGTTTGGTTGGATATACACCTTTTAGTGGTTCTTCTACTAATGAAACTTACGAGAATTTAAGATATTGGAAAAAAACTTTAAGAAGGCCCCGTAC tpg|BK006949.2|:747592-749493 7X5=94S 59=1X255=7X 
 tpg|BK006949.2| 344001 + tpg|BK006949.2| 343884 - INS TAATAAGTTGACAAATCTTCTCAATATCCCTGTCAACTGCAAAGAAAAACGACGCCAATAACTTTTGGATTTTTGGAGAGTCCAAATAATTTTGAGCACTATTAGATGAATCTCTCATTTTTGTTGGTGGCCTGCCTTCATCATAGCTATTCTTGTTATGTGCCCTATATATGTC tpg|BK006949.2|:343520-344365 7X7=80S 85S3=7X 
 tpg|BK006949.2| 271912 + tpg|BK006949.2| 272014 - INS GGCATATGCTCCTGTATGGAAAAGAGAGAATCGTAGTTTTTCGAGAGCTGTTGATACTTTGGATACTTTTTTCCAAACATCTTATCAAACTCTAACTGAGGTACACCTGTATCGGTTTGTGTTTTATATAGCATTCCAGCGTACAGTACTTGGGCAGGAGGTAGATCATGCTTTGAAACACAGCAACACAACGCTTTCAATGAGCATTCCTTCAAAGCCCAAACTCCCGCTATATATTCATG tpg|BK006949.2|:271414-272512 23S105= 37=91S 
 tpg|BK006949.2| 544209 + tpg|BK006949.2| 543988 - INS GTCTAATCATTTAGTCAAGATATTCTCTTCCCATCACTAACATCAAGAGCGCCACTTTTTGGCAATTAAACTAGACTTCTGGATGGCGCTAGCCCATTACCTACAGTACTAAAGATTATTTGCGATATTCTGATAAAGAGCCTTGAACTTCTCGGGTGACCCCCTTAGCGTTTATATAGCGGGAGTGCCAAACGAGAGGAACATCAACAACCAGTATAACAA tpg|BK006949.2|:543530-544667 7X195= 209=7X 
 tpg|BK006949.2| 492967 + tpg|BK006949.2| 493162 - INS TTCTCTCAACAATGACTGGCGACGGTAGTGCACATATTTCTAAAAACAATCAAAATCAACACAAAGATCGCTTCAAGTTTATTGTGAATGATAAAAGTATTCTAGGACCTCAATGGTTAAGCCTTTACCAAACGGATGGGAAAGTAACATTCGCAAAGTCCCACTTCGAGCAAGCAATGATGAACGTTATTAGAGAACCAAATATTAACTCTACTG tpg|BK006949.2|:492521-493608 7X77=31S 1S1=16S 
 tpg|BK006949.2| 611134 + tpg|BK006949.2| 611869 - INS TATCATTCGAGTCAACCAAGCAGCAGTTTACGCGTGTCAAAAAAATGCTGTTTCCGTTGATATGTCCCACTTCGAGTGGGCTAAGGATAAGATATTGATGGGTGCTGAGAGAAAGACTATGGTCTTAACAGATGCAGCCAGAAAGGCCACTGCTTTCCACGAGGCTGGACATGCCATTATGGCCAAATACACCAATGGTGCTACCCCGCTATACAAGGCCACGATATTGCCTAGAGGTAGGGCATTGGGTATTACTTTTCAATTGCCAGAAATGGATAAGGTCGACATCACCAAAAGGGAGTGTCAAGCCAGACTGGACGTGTGC tpg|BK006949.2|:610470-612533 7X358= 305=7X 
 tpg|BK006949.2| 284384 + tpg|BK006949.2| 284650 - INS GTGGTGTTATGGATAAGAATGAAGAATGAGGCTTTAGCCATTCATGTTTCTTGATCTGTTTCAGGTTTATTCTTTTCTTTGGGTCTGAGACCAGCATGCGTCTTAATAAGTCCCGAGGTATAGGAAGAATATAATCAGGGAACTTTAATGGTGTGGAGTTAATATAATTATAAAGTCTTCCTATATCGCTGCCTTCAGGATTATTTGGATCATCATCCCACGGTAAATATCCAGCTAGTATAGCGT tpg|BK006949.2|:283878-285156 9S66=55S 118S5=7X 
 tpg|BK006949.2| 675598 + tpg|BK006949.2| 676192 - INS GTTCTAAACCATAGAGTGGTAGCCATAAGAGCCGGCATATTGGTAATTTTCAGTATTAACGTTAGAACGTGGTGAATACGATGTGGTCCAGCCTTGCCTCGTTGTGTCATATACGATCTTTTTCTTTGGGTCACAAAGAATATCATATGCTTGAGAGATGACTTTAAATCTATGTAGTTTTTCGCTTGATGTTAGCAGCAGCGGTGATTTACTATCACTGTTGGTAACCTTTTCTG tpg|BK006949.2|:675112-676678 121S124= 222=7X 
 tpg|BK006949.2| 356121 + tpg|BK006949.2| 356888 - INS ACTTTAGACAGTATCTCATGCTACCAATTGAAAATGACGAACAAGCTAATTCAAATTGGTTTGAGAATTTTCATGCAATTGCCACGTTTGAAAACCCACATCTAATAACCAAATTTCTGAAACTGAAAAAAGGTGACATTGTATGCGGTTGTACGAGAGAGCCAAACCATTCCATTTTCGAGAATCCTACTCCCCTGGGA tpg|BK006949.2|:355707-357302 7X6=205S 175=7X 
 tpg|BK006949.2| 704306 + tpg|BK006949.2| 704686 - INS CTCACATAGTTACTATTTCTATCCGATGATCGAATTTGGTATGTAAGTTCTGTTTTTCCACTTTGCGAAGCGGTCATTGGCCCAAAAGAAATACAACGAGTCATCTCCTCACAGTAAACTGTACAACAGCAAAGAAACAGTTAAAAACCCTCCAGAGAGAACACTTACTACTATAGCATGGATGAAAACGGTACAGTAAAGCC tpg|BK006949.2|:703886-705106 7X164= 98=1X92=7X 
 tpg|BK006949.2| 109334 + tpg|BK006949.2| 109667 - INS TCTCTACTTCTTTCTCTAGAAAAAAGGCCAGAACCTTCGATTCTTCCTGGAACTGGGCTAAACAATCTTTATTATCATTATACTTTGAGATAATTCATGGTGTCTTGAAAAACGTTGATAGAGAGGTTGTTAGTGAAGCTATCAATATCATGAACAGATCTAACGATGCTTTGATTAAATTCATGGAATACCATATCTCTAACAC tpg|BK006949.2|:108910-110091 12S158= 103=7X 
 tpg|BK006949.2| 466830 + tpg|BK006949.2| 467476 - INS TGTTCTTTCGAGGACGAAATCAAATTATACGGCCCAGATGGTTTGTATGTAACATTTTGGTACCCTTTTACTGTAACTAACCTAAGGGCAGAGGTTGATGGGTTGAAGGTTATTACCACTGAAAAGATTTACTTTCTATCCAGGGTACAACCTCAGACTTCTAATATATTTAGAATTGGCTCAACCGAGC tpg|BK006949.2|:466436-467870 7X6=89S 91S4=7X 
 tpg|BK006949.2| 878574 + tpg|BK006949.2| 878218 - INS GGGAATGGAAATTAGAAATCATGGCATCATCGCCACAATTGGAAGAGGAAGCAGCTGGGAAATTAGAAACAATCCACGCATCAGCTATGGCAAAGAGCAAAAAAAAAACAGATGTTGTCGATTCAACAAACCTGCCCATTCTAGAATTACTATCATTAAAAGCTCCCATTTTCCAGTCTCTTTTACATCCTGAACTGCCC tpg|BK006949.2|:877804-878988 7X161= 188=7X 
 tpg|BK006949.2| 599983 + tpg|BK006949.2| 600259 - INS GGGATATAAACTACAGTGAAATTGATCTCAGGATCATTAGTAATTTTTCTCACTATAAGAAAAAAAAAAAAACATATATTTTGCTATGAATTATAATAAGTAAATATATACATATATATGTACAGAGAAACTGACGAAGAAAATAAATCACCCGTTAATGCTTCTTAGG tpg|BK006949.2|:599631-600611 14S103=16S 39S4=7X 
 tpg|BK006949.2| 682720 + tpg|BK006949.2| 683009 - INS CCAAGTCAAGTACGTATAAAATCTACTCATTAGTAAATCGTTGTACCCACCCCCTCCAAGTAGGAATATGTGCGCTCGAGGATAACTTTTCATGATATTTATGATGATTCGAGAAAGCCCTCGTATTGTTAGCTGCCATTCATTGAATCTATCACCCAGAAGCCCATCACC tpg|BK006949.2|:682364-683365 7X85= 183S4=7X 
 tpg|BK006949.2| 481335 + tpg|BK006949.2| 481140 - INS GCGCACAGCTCTTTAGATATGCTAAAAAAAATGAAAAAAAATGGAACAAAATATGTGTTTTTTTATTTAACGTTAAAATTAAAGATTAAGTTATTTATTCGACGTCAGCATCAAAAGTTTGACCTTCAACTAACTCTGGAATAGCTTCATCCTTCTTTTCAGCATCAGCTGGAGCCTTGGCTTCGTGCTTTTCCATTTGGGCAGCCAATTGAGACAAGGCTTGGAT tpg|BK006949.2|:480674-481801 7X5=189S 212=7X 
 tpg|BK006949.2| 366061 + tpg|BK006949.2| 366423 - INS GGCTAAAGAAGTGATATTATATCATTTTATGCACTGACTTGTAAATAAGATTATAAACGATTATTCATCTTTACTACTTGCGAACATTTCACTGTCACACCAGGCTATGAGGGCCCACAGCCAGAGAGTCGCAGGGCATAGCAGTAATACACACCAGTAGTGCAGGAAAGAGTCATTGTTGCGTAACCAGTAAAATGTAGCAAGACTAATTAGGAGTAC tpg|BK006949.2|:365609-366875 7X5=155S 206=7X 
 tpg|BK006949.2| 28368 + tpg|BK006949.2| 28890 - INS GCTTAGGAAAGTCCTATTTCATATTATTTCGTTGCCTTGTGTAAGTTAGAAGTACTTCTTGTCGATTGTGAATTCGGATAGCCGCTAGAACGCCAATCATTGCGGAGGTTTGCCATCGCATGGATACCATAGCCATCTGCACATTCTAATATAGATTATATTACTTTAGACCATGTCATTTCATAATCGTTGGTTTAAGCGGTGTTGTTTCCACAGTTTGTATGAGAACTTTTGTCCAAAGTAAAGTATCAGTAACGTAATCTGAGCAAACC tpg|BK006949.2|:27810-29448 7X158= 3S252=7X 
 tpg|BK006949.2| 33647 + tpg|BK006949.2| 34052 - INS TGGCTTTGAAAGGTAAAAAGCTTGGTAAAGCGTTACTGCAGAAGATGAATATTAAACCTGCAACAAGCCCAAATTCATCAAATGCGATTAATCCATTTTTTGATCCGGAGTCGCCAAACAAAGGAAAACTGATACTAAGTAGTGTTCCTCCCTTACCT tpg|BK006949.2|:33317-34382 7X6=73S 74S5=7X 
 tpg|BK006949.2| 800614 + tpg|BK006949.2| 801295 - INS GAGAGTACACAAAGCTATATTAAATAAAAAGAACGAAATTGGAGCTGACACCGAAGCGGAAGAAGGGGAAGAAGACAAAGAAATACAGATTCCTGTTTCTATGGCGGCGGAAGAAGAGTATCTGCGCAGCAAGGTTTTGTCAGAGCTGTTGACAGATACACTCGAAAATGACGGTGAAATGTACGGCAACGAAAATGAGGTATTGGCAGCATTGAACGGTGCATATGATAAGGCTTTGTTACGTTTATTTGCGTCTGCATGCTCAGACCAAAAT tpg|BK006949.2|:800052-801857 15S129= 127=17S 
 tpg|BK006949.2| 184257 + tpg|BK006949.2| 184288 - INS AGGATATACGATAAAAACAAGTGAACAGCTCTTACATAACAACGCACTCACTTTTCTCTTTTTCAGAAGCTTTTGCATTGAGAAGGCTGCTTCTTCGCTTAAACTTGTCTTTTTTGACTGGTGCGTGTATTTCTGAGTTTTTTTTGTGAGAATGGATTTTCCTTTTTGCTTCAAATTT tpg|BK006949.2|:183887-184658 7X4=85S 84S5=7X 
 tpg|BK006949.2| 601679 + tpg|BK006949.2| 601143 - INS AGTAGGTATACTACCAGCAATGGCACCGGCAGTTAAAAGCTCCCATGTTTTTAATCGATTCCTCTTTGTTTTATCATTTGGATCAAAATCAAAGAGATCTTTTTTTAAATGTGCATAAGTGGGAAAATAAATAGCAGAGAATGGAACATCTCTCATTAAACATGCGGCTACACCATTGTACAAGCCCCTCAGTCCTAATTTTTTGACTATTTGAGTGGCAGTTTCATTGGCTTGTTGTATGTTTTCACCAACATAGTCGGATTGGACC tpg|BK006949.2|:600593-602229 7X4=417S 252=7X 
 tpg|BK006949.2| 303806 + tpg|BK006949.2| 304510 - INS CCCTATAGTGTTAATACTTACGATGGAAACCTTATCAATGCAAGTACAACTGAATCAACGACTACTATTCGGCCTTTCGTGACTTCTCACTCCTACGTTGCTTCTTCTACACCTTATTCGAATATTTCATCATTGAATGAGGACTACGATAATGCGAGCAACTTTTTGACTCCTACAACAG tpg|BK006949.2|:303430-304886 15S51=31S 86S5=7X 
 tpg|BK006949.2| 212163 + tpg|BK006949.2| 212638 - INS TTTTTACGGCGTGTAACGGGGGCATGAGCAAATCTCTTGGATAATTCATAATCCGTGGAGCAGGTTGACGTAGCATCGTACATAGTATTATTTGTGGCAGATAATGTGTTATGATATGCTGAGACGTTTTGAACTCGTTCCACTGGGGTATTATTCGCGTTGTCATTAGGAATTGAGTTTACCAGGGTATAGT tpg|BK006949.2|:211763-213038 7X6=90S 91S6=7X 
 tpg|BK006949.2| 145799 + tpg|BK006949.2| 146356 - INS TTGAAACATATAGAATTTCATGATAATTAATTCAAACGGTATCTTAATGAGGCCAACTATTCCGGCATTCATAGACAAAAAAATTATATCAGAAACTCCAGAAAAGCTCCTACTCTCTCATCATCAATGGGCTTTCTTCAACGATATAGAAGATATACATATGTTAGTAGATAGGTTGGATGATTTAAGAGAAAATGAGGGACAATTGAAGAAAGCTTTGACATCCAAAATGGACCGTATTGAAG tpg|BK006949.2|:145295-146860 7X142= 230=7X 
 tpg|BK006949.2| 643432 + tpg|BK006949.2| 643545 - INS CGTTTCCATACTTGGTTATTGTATATGACTGTTTTCCTGATAAAAGAATGCCTGCAATAATTCAAAGACAAGAGATATAAAAGTGCACTGGCGATTTCAGGAACAATGGGCGCAACCAAAATTTTAATGGACAGTACTCATTTCAATGAGATCCGTAGTATAATCCGTTCGAGGTCAGTGGCATGGGACGCCTTAGCCAGATCTGAGGAATTGAGCGAAATTGATGCGTCTACTGCAAAAGCGTTAGAATCCATTCTGGTGAAGAAGAACATTGGTGACGGTTTATCATCTTCGAAC tpg|BK006949.2|:642824-644153 7X172= 279=7X 
 tpg|BK006949.2| 231529 + tpg|BK006949.2| 231877 - INS GCTGTTGAGCCATCATATTGATATTTCCAACATTGTGAAATCCGCTCATTTTTTTTGCTGCTATTAGCGATGCAGAATTTTTAACGATTTATTTTACTCTTCCTTCTTAGAGTAAGTATGTCTTCAACAGTCTGTTACTATTTTTTTTTCTACATACTCAATTCAGCTCTTACTGAAATTTTCT tpg|BK006949.2|:231147-232259 7X4=88S 86S6=7X 
 tpg|BK006949.2| 936050 + tpg|BK006949.2| 936443 - INS TGTGGATATGTGTTACTTTCTTTCAACTAGTTTATCGATACTTTTCGGGCTTACAGCTCCTATGTGGATATGTGAATACTCATGCTGACACTGAAGGATTATTGGTATTGGCCGGTTGTGTTTTTTCTATACATAGCAATAGTTCAAATGTCAATGACCAAAAGAATAGGAATTTTTTTAAAATACAAGGCTGATGAAGTA tpg|BK006949.2|:935634-936859 7X5=21S 176=7X 
 tpg|BK006949.2| 737529 + tpg|BK006949.2| 738111 - INS ATGGACCAATTTTGAAGTATTTGAGAAAATTCCATTATCAATAATGCCAAGTCATGAATGGATATAATTGAGCTCTTTTCCGTTTCTCCGTCTGTTTCGATATCCGACTGATTACTGTCTATATTCACATCTTCATTCTTTTGTGAATGTTCCCATTCATTTATATCATGTATAGTCC tpg|BK006949.2|:737159-738481 7X72=17S 9S1=142S 
 tpg|BK006949.2| 79482 + tpg|BK006949.2| 78763 - INS GGGTATAACTTATAGAAATGTCGTTCGCATTTGCAGCTGTCGTAGTACCAGATTCGTCATCGAGAAATTTACTCGAGGATGATTTCTCACCTCCAGAATTTTTTCCAGTTACTTCCCTATTTTCTGGACTACTAACAACCTCTTTCGTATCAGCGTAAACCTTCTCATTCTCTTTGACTGCATCATATTC tpg|BK006949.2|:78369-79876 7X5=192S 95=7X 
 tpg|BK006949.2| 914440 + tpg|BK006949.2| 915108 - INS GTGGTCGTATAGATGTTCCTTGGATTTATATTCGCAAGGGTTCTTGCTCAAATCAGTTTCAATTGCAAAGGACACTATTGAACGGATCAAGATAATTA tpg|BK006949.2|:914230-915318 7X134= 74=7X 
 tpg|BK006949.2| 74587 + tpg|BK006949.2| 74485 - INS GAGTAAGTTGCTGTCCGTCTTATCTTTAGTGTGCGTGCATTCTGACTCATCGACAATCGGGTACGATAGCGGAAAAGTTAGCAATTCTTGCTGGTAAGATTGAGAAAAGTCATCGGCATAAGTCGATCTGTCCGGGCTATGCGAGAGCATAGGGGGCTCGAAAGCAACGTTTGAAAACGAAAGAGGGAAGACCTCGTCTTCATAGCGCGAGATGGGGGAAGATTCCACAGAGGACATTGTAAATAATTGTAATTGTATATTATTGTG tpg|BK006949.2|:73937-75135 7X7=284S 134=7X 
 tpg|BK006949.2| 521433 + tpg|BK006949.2| 521544 - INS TAATAATACTACTTCAAGCTCAACAACAGCTATATGGCGGTAACAATAATAATAATAGCACCGGAATTGCGAACGATAATGTAATAACACCCCATTTTATCACCAATGTTCAATCCATCAGTCAAAATTCCTCATCTTCTACTCCGAACACAAACTCTAACTCTACTCCGAATGCAAATCAACAATTTTTGCCATTCAATAACAGTGCTTCCAATAATGGTAATTTGACGTCTAACC tpg|BK006949.2|:520945-522032 7X163= 223=7X 
 tpg|BK006949.2| 69517 + tpg|BK006949.2| 69135 - INS TTATATTCCCGCCCATTTTTTCTTCATTATCAGGTTGCGATTTTGAACAAAAAAAGTGAAACTTGAAGTTACGATGTGACATAAATTTGTTAAAATAAAAAAGATAAAATTCAGGATAGAAGTAGGTGCAACGCGAAATTGTCTCTGTCTACTTGTGCCTTGAACATCGAACTTACAACAGATTAACAA tpg|BK006949.2|:68743-69909 7X3=186S 95=7X 
 tpg|BK006949.2| 83381 + tpg|BK006949.2| 83487 - INS GATAAACCACATCCGTACATCGGCGATCGACTTGCATAGTACGTGGCACTTAGGTCACAGCCACTATTCCTTTTGCTGTTACCGCCATTGGTAGTGTTGCCAGACATTCCAAAGGGAGATGGGCCTCTACCTTGATCTTGTGCCGCCGAGGAAGGCCCATTAGTACCACTCAAGTAATTGTTCTTGTTATATGGCTGCCGCTGCGATGAGCCAAACGATATTGAGC tpg|BK006949.2|:82915-83953 7X13=100S 108S5=7X 
 tpg|BK006949.2| 165893 + tpg|BK006949.2| 165974 - INS GATTTACAGCCTCTGAGAAGACAGCATCAATTCGTATTTTCGATAATTAACTTGCCTTATAGTGTCTGATTAGGAAACAATCACGAGACGATAACGACGGAATACCAAGGAAGTTTGTGCAAATATACAGCCGGCACAAACAGCAGCTTCACTCAGGTTAACTCACATACTGTTGAAAATTGTCGGTATGGAATTCGTTGCAGAAAGGGCTCAGCCAGTTGGTCAAACAATCCAGCAGCAAAATGTTAATACTTACGGGCAAGGCGTCCTACAAC tpg|BK006949.2|:165329-166538 7X247= 258=7X 
 tpg|BK006949.2| 733692 + tpg|BK006949.2| 734030 - INS AATCATGACGTAGGTGAACTATTTTGGAAGGTCAAGGAAGAGGAAGGATCTTTCAACAACGTTATTGGCTAAATAGAAGCATCAAACATATGTATATGCACATCTATATTAATGATACATTATTCTCTTCAAGGATCCAATATGGCTTCCCATAGAATTATGAAGGAAGTCCAGTTCTCA tpg|BK006949.2|:733318-734404 7X9=81S 85S5=7X 
 tpg|BK006949.2| 933873 + tpg|BK006949.2| 933859 - INS GCTCATCTGTTATTGTATTTGAAATAGGGTCTTTGATTTCTGCTCTTTCGAATTCAATGGCGACTCTGATTAGCGGAAGAGTCGTTGCTGGGTTTGGAGGAAGTGGAATTGAATCACTTGCTTTTGTAGTTGGAACATCCATTGTCCGAGAAAACCATAGAGGAATTA tpg|BK006949.2|:933509-934223 7X11=73S 79S5=7X 
 tpg|BK006949.2| 215332 + tpg|BK006949.2| 215616 - INS CCCGCACTTCTTAACCTCTAAGGTATTCAAGGGGCGGAGGTGTAATA tpg|BK006949.2|:215224-215724 11S19= 24=7X 
 tpg|BK006949.2| 456169 + tpg|BK006949.2| 456255 - INS CCTCTTATCCCATGCTAGATCAGCTTCTTTCTCTACCTACACGTCTCCTCCTCTGTCTGCACAAACGGAATTCTCTCACTCTGCTTCGAATGCAAACTACTTTTCCTCGCAATACCTAATGTATTCGCCTCAGAAAAGTCCAGAGGCCCTATATACTGAATTCTTTTCTCCCCCTTCGTCTTCTTCTTCGTACATCAACTATAGCTATAATAACTCCAACAT tpg|BK006949.2|:455711-456713 7X154= 111=7X 
 tpg|BK006949.2| 545973 + tpg|BK006949.2| 546218 - INS GGTTTATGCTTGCGATGATGCTCAATATAAATGTGCGTGTTCTGATTGTCAAGAGTCTTGCCCCCATTTAAAACCTTTAAAAGATGGCGTGTGTAAAGTTGGCCCTCTGCCATGTTTTTCCCTTTCTGTTCTGATCTTTTACACAATCTGTGCACTTTTTGCATTTATGTGGT tpg|BK006949.2|:545613-546578 7X6=80S 82S5=7X 
 tpg|BK006949.2| 906306 + tpg|BK006949.2| 906971 - INS AGTTGCCACCCTTAGTGGTAGAGACATATTTGGATTTAAGACAGTTAAACTCGTCTCATTTAGTTAGATTAAAGGACCACGAAGGCCATTTGTGGAACGTTTGCAAAGGAACTAAGAAGCAGGAAATCGTGATGGAACGTTGGCTTATCGAATTAGAT tpg|BK006949.2|:905976-907301 7X4=75S 73S6=7X 
 tpg|BK006949.2| 564139 + tpg|BK006949.2| 563674 - INS GCTTTACACCGAATTAGATGCTGTATTCTCATCAGTTAGTTCTTGTGGCACCTATAGC tpg|BK006949.2|:563544-564269 7X13=16S 2S11=23S 
 tpg|BK006949.2| 754423 + tpg|BK006949.2| 753926 - INS CAAGTCGTTCTTGATGTTCG tpg|BK006949.2|:753872-754477 7X3=7S 10=7X 
 tpg|BK006949.2| 682067 + tpg|BK006949.2| 682266 - INS AACACAACTTTACGCCAGTTTCCCCTAACATGTTTTTTATTTCATAGCAAAGCATTTTACTCGGATCTGGTCACTAAGGAGCCGTTGATCACACCGAAAAGAATAATAAATAAGACGCCTGGGTTAAACTTATCTATTTCTGAGAGGGCTTCCAACAGACTAGCTG tpg|BK006949.2|:681721-682612 7X4=119S 83=7X 
 tpg|BK006949.2| 722019 + tpg|BK006949.2| 722434 - INS TCTATTGCCGTAGCA tpg|BK006949.2|:721975-722478 7X4=3S 4S4=7X 
 tpg|BK006949.2| 578879 + tpg|BK006949.2| 579327 - INS ATCCTTATACACCAGTTGATAAAAAGTATTGCATTTTTGAACCAATGTTTTCATTAACCCTCATTAAAAC tpg|BK006949.2|:578725-579481 7X5=30S 31S4=7X 
 tpg|BK006949.2| 929409 + tpg|BK006949.2| 929618 - INS GGCATCAATGTACAAAACACAGTAAAATCGAAGATAAGAGATGTAAAACCATAGAGACAATTTGAAAACCTATAAACACACGTTTTATACTTTATCGTTATTACGAAAAATCAATTTTTGCTCGACCAAAAGCAGCCTTCGGACTGATATATCTAGGTCCGTTAGTTTAGTAGCTGTTGAGGTC tpg|BK006949.2|:929027-930000 7X60= 92=7X 
 tpg|BK006949.2| 529368 + tpg|BK006949.2| 529801 - INS GGTCACTGGAGAATCAAAAGCATATTGCTATAATATTAACTGCCGTTGAGGAAAATATTGCAGGTCAAGCTACAAA tpg|BK006949.2|:529202-529967 11S17= 38=7X 
 tpg|BK006949.2| 540652 + tpg|BK006949.2| 540926 - INS ACCTTTTGAGTCACTAAA tpg|BK006949.2|:540602-540976 7X3=6S 2S7=7X 
 tpg|BK006949.2| 759595 + tpg|BK006949.2| 759835 - INS AAAAATTTCATTTGGATACTTTTTTGGTACGTCAATAAGACGAGCGTTTATCTTAACTGATTTTGCTCAAATATATATTGGCAAGATAACCGTGCGAATAGGTTGGAAACCCGGAATTGTGTTTCATAATGTTGATTTGAAGTTATTTGGGAAGGACAGCCATATCAC tpg|BK006949.2|:759245-760185 7X24=60S 1=13S 
 tpg|BK006949.2| 721464 + tpg|BK006949.2| 720923 - INS CATTACTGGATAGACATTACGAGAAAAAGAAAAAGGTATAACACATACATATAGAATATGTAAAAATATATAAATAAATAACATGCATTTATAACCCATGGTACTATTTTCTTCCCCTTATTCGTTACTATATTCGTCGTAACTACTGTCGCT tpg|BK006949.2|:720603-721784 11S14=1X57= 77=7X 
 tpg|BK006948.2| 798523 + tpg|BK006948.2| 798547 - INS CTGTAACTCTAAGTGCAGCTATAAATCATTTTCTTTGCTCACAAATGATTGAGGTGTTGTGCTTATACTTGCACCCGTTAGAGAGTTACAGTTTATTATGCTTATTTAATTTATTTGCTTTATATAGTTATTGTCAAGTCATCTGAACATCCCTATCCTCTTCAACACTAAGAGATTCCAAAAGCTCATCTGTCTTCTTCCTTACAAATGGGAATTCTAGAATGGTTGATAGGTTACAGCTGATCAAGCACTCTGCCTCCATACTCTTCCCTACCTGAATCAAAACTTCACATAATTTAAGCAATAATATTACAC tpg|BK006948.2|:797879-799191 7X12=171S 158=7X 
 tpg|BK006948.2| 870640 + tpg|BK006948.2| 871322 - INS AGTGAACTAAGGAGATCGATTTAGCTGTAAAGAAATACTGGATCAAATTATTTAAGAAGACTCTTTTTAAAGCATCAGAGGATTATTTTGTCTCCCTTCTGCAGGATATGCTAAAGGCTAACGCAATAGAAATTCAAAACGTTCAGAATCTCGTAGAAACAATTATAGAAGCCATAAAAGCGATTCAAAAACGTTACAATAAACCTTTATTGGACGAAATATCTCTGCCTAGACAATGCGCAGTATTTCTATGTGAAGTATACGGTTCGGATTCTTTAAATCTAATAAAAACCGCTGAAAAGAGTACCATGAAAATGACTGGACAAAAGTTGGGTCCAATAGATGCGCTAGATATGTATGA tpg|BK006948.2|:869904-872058 7X6=5S 10S340=1X6S 
 tpg|BK006948.2| 528201 + tpg|BK006948.2| 528815 - INS GGGCTAACCTGGCGTTAATAAGCCCATTGGTGAATACTTATGGGCAAGGTGGAAGAGAATCTCTACTATCCATAAATCCTCAGTAGGCTTTCCCCTAATTACCTTCATTTTTCTACCTCAATAACATATTACTCCTTTTCAATACATTTTATGGTGGTGAACACGATATATATCGCAAGGCATGGATACAGATCCAACTGGCTTCCGGAGGGTCCATATCCTGACCCACTTACAGGAATTGATAGCGATGTTCCTTTAGCAGAACACGGAGTCCAGCAAGCCAAAGAG tpg|BK006948.2|:527611-529405 25S243= 7S263=7X 
 tpg|BK006948.2| 764526 + tpg|BK006948.2| 764981 - INS TTCCTTATAAGTCGAAAGATGAAAAGAAAGAACAAATCGTATTTATGAGAAATACGCTTTGGGCCTCATTGTATGCATTTGTTAGGGACTCTCACAATTTAGTTAGTTTAGACGTTGACTATGATCAAGTACCAGACGAAATTCAATCAAGAATTGCGTTATGCTTAATGCATAATATGAAGAGAATTATGGACTCTAGCTTTAAATTAGATGAATTGACTGTACAAGATGATTTAATATTTGATGGTTCCTTGATAACTGAGACAGCAGAAGAAGTTTTGAAAAGATTAAATGACAAATCTTTACTTCAAAATGATGTTGGGAAGAAATATCTTTTAAAGAAATATTTTGAGAAAATGGAAAAGGTACATCATAATGTTCAAAAT tpg|BK006948.2|:763740-765767 7X294= 193=7X 
 tpg|BK006948.2| 218423 + tpg|BK006948.2| 218552 - INS GCCCATTACTACAGTTATTATAATTTTCTATTCTCTTTTTCTTTAAGAATCTATCATTAACGTTAATTTCTATATATACATAACTACCATTATACACGCTATTATCGTTTACATATCACATCACCGTTAATGAAAGATACGACACCCTGTACACTAACACAATTAAATAATCGCCATAACCTTTTCTGTTATCTATAGCCCTTAAAGCTGTTTCTTCGAGCTTTTTCACTGCAGTAATTCTCCACATGGGCCCAGCCACTGAGATAAGAACGCTATGTTAGTCACTACTGACGGCTCTCCAGTCATTTATGTGATTTTTTAGTGACTCATGTCGCATTTGGCCCGTTTTTTTCCGCTGTCGCAACCTATTTCCATTAACGGTGCCGTATGGAAGAGTCATTTAAAGGCAGGAGAGAGAGATTACTCATCTTCATTGGATCAGATTGATGACTGCGTAGCGGCAGATAGTGTAATCTGAGCAGTTGCGAGACCCAGACTGGCACTGTCTCAATAGTATATTAATGGGCATACATTCGTACTCCCTTGTTCTTGCCCACAGTTCTCTCTCTCTTTACTTCTTGTATCTTGTCTCCCCATTGTGCAGCGATAAGGAACATTGTTCTAATATACAC tpg|BK006948.2|:217145-219830 7X320= 316=7X 
 tpg|BK006948.2| 659274 + tpg|BK006948.2| 659918 - INS AAATATCTTTTTCCAACTTCTTTTGTTTTCTAATGAATATTTCTTTAGGTTGTTTGGATTTAAAAAATTCAGTAACTTGTTTAGCATATGGTCCTCTGAATAGGAAAAATGAGAAAGCAACAATAATATGAACATAGAAATAAACAGAGCCCCATACCATTAAAGATGGCTTCAAATCAAGGATAATAAATGGTTGCAC tpg|BK006948.2|:658862-660330 7X184=2S 1S1=156S 
 tpg|BK006948.2| 430464 + tpg|BK006948.2| 430158 - INS TCCCTTACGGATTCGCTTGATTTTCAGACCTGACATGAAATTCATTAGATTTAGATTCATCTGCAACGCTACATTTTGGACGGCAAAATCGCCAGTCGCCAATGCCACCTGATTCTCTGGTCGATTCAATGCGACATGGCGATCCTCTTCGGACGCTTCTACACCCAATGAACCAGTGGTATCTTCACCACTATCCTTAATAAT tpg|BK006948.2|:429736-430886 11S156=18S 21S5=7X 
 tpg|BK006948.2| 290957 + tpg|BK006948.2| 291068 - INS TAGCGTGTTCTCTGCACTGGCCTTATTGCGGATAGGTTTCAAATCATCCTTGTTCAAGAATTTCAAGTAATTATTTTGTAATACTCTGAACTTATTACTTTCAGTTTGTATCTTTTCTGCATAGATCTTCTGTAGATTATCTAGTATAATCAGCTCTTCTCGACTTAATTGCTTACCATCCACAAATTGAGAGTTGTATATGGTCTTTAATCGTTTCATAACAGCGTAACATTTCTGCAGCATCTGAATTACTTTGAAACTTAGATCTTCAATCAGCGCCTCATCATGAC tpg|BK006948.2|:290363-291662 7X203=50S 12S1=183S 
 tpg|BK006948.2| 169251 + tpg|BK006948.2| 169257 - INS TAAGCCAACCACGCAAATTATTGACATGGGTCCTCATGAAATAGGAATAAAGGAGTACAAGGAATACCGATACTTTCCATACGCACTTGATTTAGAGGCCGGCTCCACTATCGAGATTGAAAATCAGTATGGAGAAGTGATCTTCTTGGGCAAGTATGGCTCTTCTCCAATGATTAACTTAAGGCCACCTTCAAGATTATCTGCAGAAAGTTTACAGGCATCCCAAGAGCCATTTTACTCCTTTCAAATCGATACGTTACCAGAACTGGATGACTCTAGTATCATCAGTACATCCATTTCACTCTCTTATGA tpg|BK006948.2|:168613-169895 7X276=15S 1S1=242S 
 tpg|BK006948.2| 685101 + tpg|BK006948.2| 685242 - INS GTGTTCTTATGTATATGTAAAAGATATCAAGGCGTTTTTGAATGCGTTTTTGTTGATTTGTTTACTTTCCGGCGTATTCCTACGAAAAAAGCAAAGAAAAATACAAAAAAACGAAACATTCGCAAATGATGACAACTTGAAACCGCCAAAAGTCATCGCTTGGGAATTTTGAGGCAAGAGGCTGCTTCTATAAAAGTTTTCTTTACATGGCAAAAGGGTATTCGTATTAGGATAGTAT tpg|BK006948.2|:684611-685732 7X209=14S 3S1=323S 
 tpg|BK006948.2| 280272 + tpg|BK006948.2| 280800 - INS GTCTTGGCACGTAATAGCAAAGGGGTTGCTTGAAAAAGCATTACATTTAGAATCTGAATTATTCGACAAGTCAAAGGGATTGATTTGGAAGTCTTTTTCCAATGAAGTTGAAGCCATTTTTTCGGAAAGGCTATCAACGTTTTTATTCTTCTTTACTCCTCTGATACAGCGAACAGAATTGCCCTTCCTTTGACATTCGGTACACAGGAAGAC tpg|BK006948.2|:279832-281240 141S174= 9S191=7X 
 tpg|BK006948.2| 551115 + tpg|BK006948.2| 551681 - INS TTAAATACCGGATGTGACTACATATAAAAAGTGCGCCTTTTACAGTGATAATTAGCGTCAATCAATAAAATATTTGTAAAATAGGAAGCGAAATCCCGCAGATGCCAGAATAGGTGGTGTATAAGGCAAGAAAACTTTACCTGCATAAATTAGTATTGAACACCAATCAAGTAGTCAGCCAATTGCTCGACAATCTTGGTGGCCTCACCGGCTTGTACGGTTGGTGGATAATGAGCAATAATAACGGTTTGCTTAGTTCTTACACAAACAACACCCTCAGCATCATGTCTACCG tpg|BK006948.2|:550513-552283 7X135=85S 1=187S 
 tpg|BK006948.2| 149749 + tpg|BK006948.2| 149050 - INS TCTAGCTCCTATACATTGAGTTGTCGACAGTAAAAGCTGGTATATTTTTTAGTACCAAACAATTAAAGTCAATCGCCAATGAAACCAATATTCTTCAAAAGGAGTACGACAAGCAACAATCGGCTCTGGTTAGAGAAATTATAAATATTACATTAACGTACACACCAG tpg|BK006948.2|:148700-150099 7X4=355S 147=7X 
 tpg|BK006948.2| 478713 + tpg|BK006948.2| 477995 - INS TTTCATTGCCAAGGCGATAATGTGGTCGACATTGAACATTTCAGAAAGACGAGAAATGGGCATGTCATTATCTACAGATCCGTCCATGAATTTCATGTTTGATAAATGTAAATTTGTTGCCCCCCACTCTTTAATCTTTCCAGTGTGAGGATCTTTCTCGAATAGCGGCGTGGAGGGGAAAACTCCAGGTAGAGAACAAGATGCGCATACGGCAGACCAGATGAGAACGTTTGGAGCGGTTAAATTGTTTAGTAGTTTCGGCTGTTCGTATATGGAAGCAGGCGAGACTGTGATATTCAGGATTTTTCCAGTCTTGTTGTAGGCTTCCCTAAAGGTCAAGTTTCCTAAAAACGAAAGCATTGTGTTAATCAAAGGTTGATTATTGAACCAGGTACCGTTTTGGCAGAACCTCGATATCTTGATTAGTAAGTTTTCGTTGGGAGATTTGGAATTGTCGTCATTGAAGATGTTAAACTCCATATTAAGTACATTGGTCAACAAGGAGGGAATTTCCTGGGTCGTGTGGACGCAAAATATGCTGGCAACAATGGCGCCAGCACTGCTACCGCTGATCACCTTAGGCATCAGGTC tpg|BK006948.2|:476799-479909 7X5=216S 573=7X 
 tpg|BK006948.2| 395738 + tpg|BK006948.2| 396276 - INS GCAATGAACTGTGATGTTGTTGTGGAACCTGTCCATGCAAAATGTGGGTTATACCTACTATTTCCTTAATAGTAACGAGCCATTGATTAATACCCATCATTGAAAAGCAAGCGCTAAGAATGGCGCGGCGCCTATTTCTTGGTTCCAAACCATCAA tpg|BK006948.2|:395412-396602 7X4=74S 73S5=7X 
 tpg|BK006948.2| 768875 + tpg|BK006948.2| 768978 - INS GGTTCAGCACGGGTGTCATCAAGCTATGGGATGCGCGTGCTGTGCAACTGGCTACTACTGACCTCACACATAGGCAGAACGGCGAGGAACCGATCCAAAACGAAATAGCCAAGTTGTTCCATTCTGGCGGCGATTCCGTTGTCGATATCCTGTTCTCACAAACCTCTGCAACAGAATTTGTTACGGTTGGAGGAACGGGTAATGTCTACCAC tpg|BK006948.2|:768437-769416 7X86=20S 16S1=225S 
 tpg|BK006948.2| 312923 + tpg|BK006948.2| 313199 - INS TGGCTTCATCTTCTTTCGTCAAATCGTCGATTTCTTCGAAATATTTTGGCTCTTTCTTTAAAAGATCCTTATCCAATTGTAAAATGGCCCTCTTGCAACGAATCTTTTGCCATTCCAACTCTTGTATTCTATTATTGGCCTTTTCCACTGTTTGTGCATGCCCCTTCGTGACAGTCCTTTGATGGTTACATAGGATG tpg|BK006948.2|:312515-313607 7X75=23S 10S1=265S 
 tpg|BK006948.2| 968807 + tpg|BK006948.2| 969288 - INS TTGTATCTCACCTATCTTTCAAAATATTACTATTCACTCTGCTAAGATTATCGGAATAGGGACCAACTATCATCCGCTAATTACTGACATTACCAAATGAGATCTGTGAATGGGCAAGATAAAAAACAAAAATTGAAATGTTTGACGTTATGTAAAACTATTAATTCCTTCGCTTTCGGCGGTCACAGAATTTGCGTGTAGCTGACTCTTGTTCAATCAATATCATTTGTTACTTTATTTGAAAGTCTGTATTACTGCGCCTATTGTCATCCGTACCAAAGAACGTCAAAAAGAAACAAGATAATTTTTGTGCTTACACCATTTATAGATCACTGAGCCCAGAATATCGCTGGAGCTCAGTGTAAGTGGCATGAACACAACTCTGACTGATCGCACATATTGCCGTTATCATAAATACTAGTTGTACTTGTCAATGCGACGAATGGCATCATGCCTATTATTACGTTCCTCTTTTTCCGTTTCATGTTTCCAGAATGCTATTGAATCTAAC tpg|BK006948.2|:967771-970324 7X344= 256=7X 
 tpg|BK006948.2| 868131 + tpg|BK006948.2| 868894 - INS TTATATCATGCCTTATGATAGTGAAAGACGTTGTTGCTTCCTACTTGCGTCCCCAATCGATCCGCTAACCTTTTTTTTAACTACAGCATAACCTCACATCTACGTATCCTTACATCTATAATATTTTTAAATAATTGTAAATTAGAAAAACATCAAAATTCCGTTCTATATTTTGATACATTTTGTTGCAGTAGTCCAAGATGAGATCAGAATAAGATAGGTGAAAATTTTAACAAGTACTAAAGCGTTCGTTGACAGCTTTCTTTGCGTTGCCATGGCTGAATTAAACGATTATAGTACGATGATCGATATTCTTCTCTCTGATATGGATTTGGAAACGGTCACAACTAAAAAGGTTAGGATGGCTTTGAAAGAAGTATATGCAATCGACGTTGAATCACAGGG tpg|BK006948.2|:867307-869718 7X374= 203=7X 
 tpg|BK006948.2| 286530 + tpg|BK006948.2| 285867 - INS ATTGTTGCTTCATATTTGTTTGTATATACATCTGAGCATTGCGGATCTAAATAGTGTGAAGTTTTTGAGGTGACTGACTTTCTCAACACGTCGAGCACGACATTTCCCAAAAATAGCTGAAGAACATAAGCTAAGCAAATTACGCAACACACTCTCATATGACCGAAGACTTTATTTCTTCTGTCAAGCGT tpg|BK006948.2|:285471-286926 7X5=232S 180=7X 
 tpg|BK006948.2| 364157 + tpg|BK006948.2| 364335 - INS TATTGTCAATTACACCATTCGCTTCTCTTCCTCCATAAGTAATAATGTTTTCATCATCATCTCGACCTTCAAAAGAGCCATTACTATTTGACATCAGACTTAGAAATTTGGACAATGATGTTTTACTGATAAAAGGCCCCCCTGATGAGGCATCTTCTGTCCTACTATCTGGAACTATAGTATTGTCAATTACTGAGCCAATTCAAATCAAGTCTTTGGCTTTGAGACTTTTTGGTAGGTTGAGACTAAATATTCCAACGGTTTTACAAACTGTTCATGGGC tpg|BK006948.2|:363579-364913 7X4=341S 265=7X 
 tpg|BK006948.2| 1031676 + tpg|BK006948.2| 1032451 - INS AACCTCAGTGTACGTTTCCCACGAGAAACTACAGGGATATTTATCTTCCACATGTCATTCATAGCTTCATACTTGTCGTCACCAGTCTGACTATACCCTCCAAAGATCAGAATGGTATTAACAGATGAGCAAATGTGTGTTGCTGTGCTACAATGTTTGGAAGAGAGACTATCTGTAGACCTTGGGTTTGTTACAGGTGGAATTGCATCATCCTCTAAATAGTCCGTACTTCCTGGTGAACCAACCAAATCATCTATTTTGTGATCCCCATTACCTTGGCGATATGGGCTTATCGACCTTCTTCCTTTCGCACTTGTTGTGGTATTTTCATTGGATACATTGTTGTTGGAATTACTTATTGATGCCTGCATGTGACCAAATCTTGGCGAGAAATTATTGTAAATTGCAAACTGGTACGGAGGAGCGACTAATTCAATCTTTGAGAAATTGAACGTCACTGTATCTAGAATGTAACCAGTAT tpg|BK006948.2|:1030700-1033427 7X279= 466=7X 
 tpg|BK006948.2| 920908 + tpg|BK006948.2| 921093 - INS GCACAGCAAGCTATAACGTTGCTCAACTTTTGATTCCGAAATCAGAAGCTTAAATAAGGAAAACTGAAAGCTAATTGGATGAAGCACACAAACTTAATCAACCTTATTATTCAAAGTATTCGGAGCCCTAGTAAAAACTGCCTATGATATGTATGAGTCGTGCTTTTCCGTCTGGTTTAATAAGTGTTCGAGTCAGCTCAAATCGCATTTTTGTCTTGAAGCTTCCGCCAAAAGAAAAAAAAAGTCGTTAATAGCGATACAAGTAAGCAATTAACTATCACACCATAGAATGAGTTGACAAGAGTACTTATTTGATGGCTTTACTGAACTATGTATACA tpg|BK006948.2|:920216-921785 7X8=212S 170=7X 
 tpg|BK006948.2| 141046 + tpg|BK006948.2| 141568 - INS CATACTAGCCATGAACTGGAGGCTAGTAACATTTTCTTCACTATTAGAGGGTGAGGAGAATCAACAATTTTGAAGACATTGTCTGCGTTCACTAAACCGTGTCCTGCTACTGTACTTTGTAGATTGTTTATGGCCTGTCTCATGTCACCCTCCGCTGTAAAAATGATTGCTTCTAACC tpg|BK006948.2|:140676-141938 23S73= 40=56S 
 tpg|BK006948.2| 809369 + tpg|BK006948.2| 809396 - INS GTTACTCCTTGTCTCGTGGAGATTGGGATAGTTGGAATATGAGTTTGACGCCAAAATTTATGATCCTTTTCTTCTACAGGAGAACCATCCCAATTCAATCCTGATGCATCACCAGTCGAATATTGGGGCAATCCTACAGGCTTAGATTGAACAACGTCTATATTCTCACCATATGGCTCAGATATGAAGATTACAGCTTTAGCTCCGAATTTCTCAGCAATTAGTACTTGCTGACTCACTAATTTATCATATTGCAGTAAAAGCACATAGTCCTTCCCATCTTCTATCGTTTTCGAATCTTTTAAATGTTGTAAATCGTATGGTGTACCTTTG tpg|BK006948.2|:808689-810076 7X230= 156=1X10=7X 
 tpg|BK006948.2| 255205 + tpg|BK006948.2| 255401 - INS TTGGTGTGTCGACGCTGATGGCCGGCTTCGACCCGAGAGATGATGAACCCAAGCTTTACCAGACCGAGCCAAGTGGTATATACTCTTCGTGGTCCGCTCAGACCATTGGGAGAAACTCCAAGACGGTACGTGAGTTTTTGGAGAAGAATTACGATCGCAAAGAACCACCAGCCACAGTGGAAGAATGTGTCAAACTTACTGTAAGATCTCTGTTGGAGGTAGTTCAAACAGGTGCAAAAAATATTGAAATCACTGTTGTTAAGCCGGACTCAGATATTGTTGCGTTGAGCAG tpg|BK006948.2|:254607-255999 7X19=1X253= 201S6X1S 
 tpg|BK006948.2| 373331 + tpg|BK006948.2| 373495 - INS AAATTCCAAAACTTTAGAAGTTAGTCCATAAGCTTCACTACAATGTGGTAAATAAGTTTGTTCGTAATGAGCCATTTCTTTACTAACAAGAGGTTCCATCCTATAAGAAATGGGATCACAGACGTGGTAAACATTATAAATGTCCTTACATTGCGGTCTCTGTACGGT tpg|BK006948.2|:372981-373845 7X5=79S 80S4=7X 
 tpg|BK006948.2| 846662 + tpg|BK006948.2| 846917 - INS CGTCTTCTAGTTCATCGTCTTCTAGTTCTTCCAAATCCGACAAGTCTTTATCTTCTAGTCTATTTTCATGCTGCTTGGCAATTGCTTCTTCTAATGCTTCTTCTAACTTTGCAGTGGGCGAAGGTGCACGTTCTGGTATTACACCCTTCGCTCTTAAAATATCGTTCCATTCACTGTCTTCAGATTCGTCCACCTGGACCTGAAACATTGGTTCATTCTGCATTATGTCTGCTGAATATGCCTTTCTTCTCAGTGATGTTTACTCGAAGGCGTTATCTTGTACTGCAGATTTCTTCAGGT tpg|BK006948.2|:846048-847531 7X529= 282=7X 
 tpg|BK006948.2| 867276 + tpg|BK006948.2| 867303 - INS TCCTATGATCTTTGTACTAACTTATCTTCAATTTCAACGGAGAGATGTAAACATCATTCTCTCCTATGATAATTTCTTTTTTTATACAGAAGGTGTTGTTGTCGCCAAGAAGGATTTCAACCAAGCCAAGCACGAAGAAATTGACACCAAGAACTTGTATGTCATTAAGGCTTTACAATCCTTGACTTCTAAGGGTTACGTCAAGACTCAATTCTCATGGCAATACTACTACTACACCTTGACTGAAGAAGGTGTTGAA tpg|BK006948.2|:866744-867835 7X231= 130=7X 
 tpg|BK006948.2| 1011391 + tpg|BK006948.2| 1011931 - INS GTCATGAAGACGGATGAAGATGTCAAGATGATTAGTGCAGAGGCCCCCATCATTTTCGCCAAAGCCTGTGAGATCTTTATTACAGAACTGACTATGAGAGCTTGGTGCGTGGCAGAAAGGAATAAAAGACGAACTTTGCAGAAGGCAGATATCGCAGAGGCCCTGCAAAAGAGTGACATGTTTGA tpg|BK006948.2|:1011007-1012315 7X4=88S 81S7=1X4=7X 
 tpg|BK006939.2| 116494 + tpg|BK006939.2| 116166 - INS ATATAAATCAGCATCCATGTTGGAATTTAATCGCGGCCTCGAAACGTGAGTCTTTTCCTTACCCATGGTTGTTTATGTTCGGATGTGATGTGAGAACTGTATCCTAGCAAGATTTTAAAAGGAAGTATATGAAAGAAGAACCTCAGTGGCAAATCCTAACCTTTTATATTTCTCTACAGGGGCGCGGCGTGGGGACAATTCAACGCGTCTGTGAGGGGAGCGTTTCCCTGCTCGCAGGTCTGCAGCGAGGAGCCGTAATTTTTGCTTCGCGCCGTGCGGCCATCAAAATGTATGGATGCAAATGATTATACATGGGGATGTATGGGCTAAATGTACGGGCGACAGTCACATCATGCCCCTGAGCTGCGCACGTCAAGACTGTCAAGGAGGGTATTCTGGGCCTCCATGTCTTGCGAACGTACATAACATGTCCTTTTTCGTTGTAAAAAAACAACCAAAATAAGTTTAGGACACTTTATGGGTTTTATTGGGACATTTTATGGTTTTTTTGGGACGCTTTATGATTTCAGCGACAGGTGCGATAATCCTTTCGCAAAAACTCGGTTTGACGCCTCCCATGGTATAAATAGTGGGTGGTGGACAGGTGCCTTCGCTTTTCTTTAAGCAAGAGAATTTATAAATGTGGGGCGGGCTCTAACCACATACTTAAGATGTCGAAAGCTACATATAAGGAACGTGCTGCTACTCATCCTAGTCCTGTTGCTGCCAAGCTATTTAATATCATGCACGAAAAGCAAACAAACTTGTGTGCTTCATTGGATGTTCGTACCACCAAGGAATTACTGGAGTTAGTTGAAGCATTAGGTCCCAAAATTTGTTTACTAAAAACACATGTGGATATCTTGACTGATTTTTCCATGGAGGGCACAGTTAAGCCGCTAAAGGCATTATCCGCCAAGTACAATTTTTTACTCTTCGAAGACAGAAAATTTGCTGACATTGGTAATACAGTCAAATTGCAGTACTCTGCGGGGGGTGTATACAGAATAGCAGAATGGGCAGACATTACGAATGCACACGGTGTGGTGGGCCCAGGTATTGTTAGCGGTTTGAAGCAGGCGGCGGAAGAAGTAACAAAGGAACC tpg|BK006939.2|:113942-118718 594S11=274S 119S320=3I111=7X 
 tpg|BK006939.2| 335664 + tpg|BK006939.2| 335446 - INS GGAGGGAAGAGTGTAGCTGGTCTCACCCTCTGGCCGGGCCGGTCCGTTTTTGTGGCGTCGCTGCAGGTAAACGCGCAGTTTCTGCGCGTTTACCCCTGAGGTGAATACCATCTTCAAGCGTCAAACTGCATCCGGATATCCTGCTGTTGGTAGCGATGGTGGTGGTAGTGGTGTATGCTCTTGGTTCTGGTGGTGTCTTGCGTCTTCTCTTCTCTTTCTGTTCGTTCGGTTCGTATATAGGTATGTATATATAATGAAGGATGGAAGATCCTTCATTGCAAGTGGGAACGGCCGGCCTTGTGGTCAGTGTTACTGTCATTCTCGGGATGGGAGGAAGCCGGGTCATGGCCCATGGTTTGGAGCAGTTGGGCCAAGGCAGACTGGGGAAGAGTGTAGGTG tpg|BK006939.2|:334634-336476 7X521= 375=7X 
 tpg|BK006948.2| 680595 + tpg|BK006948.2| 681089 - INS GAACTATATGTAGTAAGTGGACGGGCAAAAAAAAAAAAGCGCCAGCAGGAAGAAAAAAGGAATCTAGTAAAAAATAAAAATTAGGTTTATAAAGTAGTAAGTGAAGTGCAAGAGGGAGCGTTATTGGACGATCATATTGTGATCGGATCCCGTTTATTGGTCTTTGATTCAATTTAAAAGAAAAGAAATGTACAGGTTAAACT tpg|BK006948.2|:680175-681509 7X183= 5S186=7X 
 tpg|BK006939.2| 470305 + tpg|BK006939.2| 470733 - INS GTGTTGGAAACTTTGTTCGTCAGGTTTGACAGCATCGGCAGTGGCGCAGTGTTGGAAACTCTTGGATTTTGATGATTTTTTTGCATCACTTTCCGTGGTTTTTTCAGCATCATCAGCATTCTCTAGGAATTTTTTCTCATAGGTTTCCTTATCGAATTGCTTATACATAGTCAAACAAGCATCTAATAATTTACAGGATGATGTGCCGACTCTTGAATTGGTATTCCGTGTACTGAGAACGTTAATTACATCAATAAATGGCTTACAGTAGAGTAACACTTGTAACACAGAACTCATAAAACAAATGTTGGCTCTGTTAATTATGCCTCTTGGAATAATGGAATGGACTGGTATTTTGTTTTCAACATCTTTATTCCGTAAAACGTAACTAATGAAATCGGGATCAAAACACATTCTTAACGCAATCGAACCCAGTGGCTCAATACCCTTTGTAGAAGGTGGAACGTATTTTTTATCCTTTTTCTGAGGCTGCTTGGACAACAGGGGAGAGCTGGATTTACCTATAGTCGCCGCAGCCATGTTTGTTGATGAAACGCCTGCGGTCGTACCAGAAATTGGTGTTTTAGTGACCATCGATCCGGAGACTGTTTTGTTACTAGCTTGTCTACTTTTAATCGCATCTGATGCTATGGCGGACCAGGATTTTGCTGCTGGAGGAG tpg|BK006939.2|:468931-472107 7X586= 659=7X 
 tpg|BK006939.2| 356546 + tpg|BK006939.2| 356704 - INS CCTACAGAGTGACAATATCACCTCAAGGGACGAACCATTTTTAGACTTTCCAATAGAAGTACAGGGTGATGAAGAGACTGATATCCAGAAGATGTTAAAAAGCTATCATCAGCGTGAGATGTTGAACGGGGTTAACAAATTTTATTGTAACAAATGTTATGGTTTACAAGAAGCAGAACGTATGGTCGGACTGAAGC tpg|BK006939.2|:356138-357112 15S90= 89=17S 
 tpg|BK006948.2| 675597 + tpg|BK006948.2| 676087 - INS GCATAAGGCTCCTCCCCCTCCTCCGCCAACGGCCGAAACATTTGATTCAGACCAAACAAGTTCATTTTCCGATATCAATTCGACAACAGCATCCGCACCGACTACCCCAGCCCCTGCTCTTCCTCCTGCATCTCCTGAAGTAAGAAAAGAAGAAACGCATCCAAAGCATAGTTTACCGCCTTTACCAAATC tpg|BK006948.2|:675201-676483 7X5=90S 91S5=7X 
 tpg|BK006948.2| 693033 + tpg|BK006948.2| 693519 - INS CACAGCAAAGACTACGATTCCGAACTTGACCTACCCAATATTGACTTGAATAACTCAGTAATAAAAGAAGCAAGTGGCAGCAATTCAATTCCTACATCAGAAACAGACGCACAATCCTCGAGTTCGTCAGTTCTTCAAGGAACTATCATGACAGAACAAGCTACTCAATCCTCTCAACACGAATGTAACAGTTCACTTGATACTCTAAAAAAAAATCATCAAAAATTATTGAAGGATTTGAATTCTAGAGAGTCTGAACTACGTAATGC tpg|BK006948.2|:692481-694071 5S2X89=1X194=1X23= 7S246=7X 
 tpg|BK006948.2| 1021030 + tpg|BK006948.2| 1021704 - INS AAATGGTTCAAGGCTGGAAAGTCAGATGGGTCACGATGTAATCCGATAGACGTCCCTATTAGTATGACAAGGTTAATTATAACATCCGACGGTTGTTCTAACAGAAAATCACCCTCAGTTGGGGAAAAAACAAATGCACACCAGATATAGAGTAAGCATGAAATGGTATTTTCATTTGCACAAGCACACCAATTTTCCGATGCAAGTATCTGCTGCGCTAGGAAAATTACTTCGCTTTGAATCGGATATTGCTCTAGCATCTCTTTGGTAATATACGGACTGTAATCTTCAATCTTATCTTCTATAAATGTCAAAGAGATATACGCGATCCTCAAAATTAACAGTAAGATACACAGATTCTCCATTTTATTTCGTATAAGGGTTGTGCCCATCGAT tpg|BK006948.2|:1020224-1022510 7X305= 198=7X 
 tpg|BK006939.2| 235072 + tpg|BK006939.2| 234989 - INS CAGTTATTGAACCGTATAGGAAGAGAGTTTGTGGTGGTGACACAGATTTTGCGGAGGTTTTACAAGTATCCTATAATCCCAAAGTGATAACTTTGAGAGAATTAACTGATTTCTTTTTTAGAATCCATGATCCTACTACATCTAATTCACAAGGACCTGATAAAGGTACACAGTATCGCAGTGGATTGTTCGCTCATTCAGATGCTGATTTAAAAGAATTAGCCAAAATAAAGGAAGAATGGCAACCAAAATGGGGTAATAAGATTGCCACAGTTATTGAACCAATCAAGAACTTTTACGATGCTGAAGAATACCACCAGTTATATTTAGATAAGAATCCACAGGGATATGCATGCCCTACTCATTATCTGAGAGAAATGTAGCTTTTTTAGTGTACGTGCCCTTATTTATGAAAAAAAGTCAAGTGCATGAATGAAATATTTACTGTTGAAGAATTTATTATATATATAGGTATACAGGATCTATCTTTTCGATAACGTAACTTAGTATCACATGTATTAGTATTAATACTGTGATAGGA tpg|BK006939.2|:233893-236168 7X218= 4S521=7X 
 tpg|BK006939.2| 312876 + tpg|BK006939.2| 313072 - INS AGGACTCAGGTACAGTACCATTTGCAGTTAATCCTATCGTCTGGTAAAATTCAACCATAGAAACTGGAGCGATTGCCAAATCATCGTCCATTTGCCAGAATCCTGATGGCAAGCCCTGGCTTTCACCGCCCGTCAGGTAGATCTCAGCACGTGTGCATGCGCATAAC tpg|BK006939.2|:312528-313420 7X136=13S 1=206S 
 tpg|BK006948.2| 374870 + tpg|BK006948.2| 375327 - INS TTAGGGAATATGCAAAAAAATACAATCCACTTTTTCTTCCAAAGCGACAAATTAGGTCAGAAAACCAACAGAATATTATATTACGTAATTTACTTATTTATATGTGTGTACTATGTATGAGAACCACGCAGTCTTGATTTCGACCTTAGAT tpg|BK006948.2|:374554-375643 7X4=71S 71S5=7X 
 tpg|BK006948.2| 759841 + tpg|BK006948.2| 760057 - INS CTCCATGACCCGGAGAGGCATTACTTCGATACTGCTAATAACTCTAACGTCGCAACAGGCACCAGCGCGGCACCAGAGCAGAACAACTACTATATTCATTGTATAATTGGTACAGAGGAGCTGACACAAGCAGAGTTAGCCAACGAAGATCTAAAGGACGATGCAACTCCGTCCAATGACTCCATGACCACGCAGGCCATCGGGTTTGATAGGCTACGATCCGTGGGATTTAC tpg|BK006948.2|:759361-760537 7X193= 38=1X165=7X 
 tpg|BK006939.2| 205466 + tpg|BK006939.2| 205133 - INS GTATATCAATCTCGAACAACCATTAAACCCTGATTTTTCAAAATTAAACCCACTATCCGCCGAAATTATCAACAGGCAAGCTACAATAAACATCGGTACCATCGGTCATGTCGCCCACGGTAAATCCACAGTAGTTAGGGCTATTTCAGGTGTCCAAACAGTCCGTTTTAAGGATGAATTAGAACGTAACATTACTATTAAGTTAGGTTACGCTAATGCTAAAATTTATAAATGTCAAGAGCCTACATGTCCCGAACCTGATTGTTATAGATCATTCAAATCTGATAAAGAAATCAGTCCTAAATGTCAAAGACCAGGTTGTCCGGGGCGTTACAAATTGGTCCGTCACGTTTCTTTTGTTGACTGTCCCGGTCACGATATCTTAATGAGTACTATGTTATCAGGTGCTGCTGTTATG tpg|BK006939.2|:204283-206316 7X279= 405=7X 
 tpg|BK006948.2| 631127 + tpg|BK006948.2| 631817 - INS TGACAATACTCTTTACTATACAAACTCTCCACCTCAACTGATCACCCTTCTGCTGAATTATTAGTTTATCCTTTTCATCTTTCTTTTTGGTATTTTGCCACTCGGCCGGGTTATAAAATACGAAACATGGCCCTAATTTACCCGCTTTTACAATAAAGGGTTTGTAATGAGGGTAAAAATATTGGCCCTAATGAAAAATCACTAGCAACGGAAGTGCAAGTAGAACCCTGAAGTCGCCGAGTAGGAAAGTGATTCCCAAGAGGAGTAGAATAAAGAAGAGAATCTACATATGGATTATTTAGGTAATAGTTTCATTGCTGATTGTCAACAACAATAATAACAAGGATAATTGA tpg|BK006948.2|:630407-632537 7X353= 331=7X 
 tpg|BK006948.2| 447233 + tpg|BK006948.2| 447352 - INS GTGTAACACTATATCATATAGTGTAATGAAAATGCAAATTGTAAAATAATATTTTACAATTTGCATTTTCATTACACTATATCATCTACTATTTTTTCTCAGAAGCGGAAGTTATAACTAATTTGACAATGTTTTCAAATCTATCTAAACGTTGGGCTCAAAGGACCCTCTCGAAAAGTTTCTACTCTACCGCAACAGGTGCTGCTAGTAAATCTGGCAAGCTTACTCAAAAGCTCGTTACAGCGGGTGTTGCTGCCGCCGGTATCACCGCATCGACTTTACTCTATGCAGACTCCTTAACTGCCGAAGCTATGACCGCAGCTGAACACGGATTGCACGCCCCAGCATATGCTTGGTCCCACAATGGGCCTTTTGAAACATTTGATCATGCATCCATTAGAAGAGGTTACCAGG tpg|BK006948.2|:446391-448194 7X161= 15S372=7X 
 tpg|BK006948.2| 758594 + tpg|BK006948.2| 758644 - INS AGATAGGAGTTCTAGTTCTTCTGCATACTACTTAGTCCTCTTCTGTCGTTGACATTCAATTGCTTGTGCATTTCTAACATGAAATAGTGGTACTACGAATGCTATTATTCTATGCCAGGCAAATTCCTCTGGAACTTTTTTTTTTTCAGTTTTTTCGTGGTGAGCTTTTTTTGCCTGTCTATCTCGAAAG tpg|BK006948.2|:758200-759038 7X5=90S 90S5=7X 
 tpg|BK006948.2| 342752 + tpg|BK006948.2| 343323 - INS TTCTGAATGATTATAAAGGGCAAAGTAGCTTGCACCTTTTGCGCTACACTCACTGTTACAGTGTGAACTCGACTGCCAGTTATATGAATCGGCCTTTGAAAAGTCAGAGGGTAGTGAGCTAAAACAATTCACGTATTCATAGGCGTTCGCTTGCGATAAA tpg|BK006948.2|:342418-343657 7X5=75S 73S7=7X 
 tpg|BK006948.2| 161499 + tpg|BK006948.2| 161598 - INS GAAATATGTGCATAGGAGAAGTGCAATTGCGTAAACTCGTTTTTTCGGCGCCGCAAAGCCAAATACATCATATCAACACTTTTCACTTTATTTTTCGTTCGACCCTTATATTTGTCTTTTGCCTTCATGCTCCTTGATTTCCTATTTCATTTACCATCATTTCTTCGATCCCCCTCATCG tpg|BK006948.2|:161125-161972 27S66=4S 84S6=7X 
 tpg|BK006948.2| 754090 + tpg|BK006948.2| 754409 - INS GCTGTGGTGGGTATTAGAATAACAAGTAGAACTAAAACTGATAGTGCTATTAATGTAAAGACTAAGACATAAGATCTTTTCTCGGGCAGAGACCATTCTCCCCATCGACGATTAAATTTGTTTACACTGAAAAAGGAATGCGTGTGATGCTGGTTTTCAATATCATTAAACTGGAAGCTTTCTCGTCTGGGACGCATTGAGTATTGTTCCTGGAGAAAGGGGGTTTGAGGAACATCTGTAACATCTATTGTAGCTTCTGTCGGTCTAATCTCGTTAATTGTATGTCCATTCTCGTTACTTTGAGGATCTGTGTTAGCTACACTATCGTTATTAGGAAAGAATGGCTTATCCATGGAAGAGGTTGAAC tpg|BK006948.2|:753342-755157 7X167=1X28= 338=1X6=7X 
 tpg|BK006948.2| 964966 + tpg|BK006948.2| 965118 - INS TTGGAAGACAGATGTTATCCATAGACAGATTCCTCATATTGACCGTTGTGTTCATCCAGAACCTGAAAACGGAAAACGTGTCCTTGTCACAGAAGGTGTTAATTTCCAAGCTATGTGGGATCAAGAGGCATTTATCGACGTTGATGGTATTACATCTAATGATGTTGCTGCTGTGTTGAAAACGTACGGTGTAGAAG tpg|BK006948.2|:964558-965526 28S47=30S 93S6=7X 
 tpg|BK006948.2| 649329 + tpg|BK006948.2| 650025 - INS CTTAAAGGAACACCTTGAGGTTACTGGTGGCAAAGTTCGTACAAGGTTCCCTCCGGAGCCCAATGGATATTTGCATATTGGTCATTCTAAAGCTATTATGGTTAATTTTGGCTATGCTAAATATCACAATGGTACCTGTTATTTAAGATTTGACGATACCAACCCCGAAAAGGAAGCTCCTGAATATTTTGAATCCATTAAGAGAATGGTTTCTTGGTTAGGTTTTAAACCATGGAAAATTACTTACTCAAGTGATTATTTTGACGAGCTTTATCGCCTCGCTGAAGTGTTGATCAAAAACGGCAAAGCTTACGTTTGTCATTGTACCGCCGAAGAAATTAAAAGAGGTCGTGGTATTAAAGAAGACGGTACTCCAGGTGGGGAGA tpg|BK006948.2|:648543-650811 7X238= 193=7X 
 tpg|BK006939.2| 277311 + tpg|BK006939.2| 277333 - INS GCTCTGGGCGGGTAGGGGGTGCAACTACTGCAGGTGGTGTTCTTTCTTTTGGTTCATCTGTTTTTGGGTCAGCTGCGGGTTGGGCGACTTATGCAGCAGATTACACTGTTTATATGCCAAAGACCACAAGTAAATACAAAATTTTTTTTTCCGTAGTAGCCGGTCTAGCGTTCCCTCTATTTTTCACCATGATTCTTGGTGCTGCTTGCGGTATGGCGGCCCTTAATGACCCAACCTGGAAGTCATATTATGATAAAAACGCCATGGGTGGTGTCATATATGCTATCCTGGTCCCTAACTCTCTAAACGGATTCGGTCAATTCTGCTGTGTTTTGTTGGCTCTTTCAACTGTTGCTAATAATGTCCCTGGAATGTACAC tpg|BK006939.2|:276539-278105 7X7=183S 356=7X 
 tpg|BK006948.2| 240314 + tpg|BK006948.2| 241038 - INS TTTCTTACAGTATAAATGCTCTTGAGTTGAAAATTTCTTTAATGAAGTTTTTTCTAAGCAGTTCGTATCTCACTTTCATTGTTGGTATCGTTTCAGGAAACCAAATATCAAACTGTCTTATGAAAATCTTTAGCCAACGACTTACGTTACTTTCCTTTGAAGAACTGTGTTCTTTGAATTGTCTTTTTAAACGTTGTGGCCCCTTTTCTGCAAGGGTCATAGAATTAGCA tpg|BK006948.2|:239840-241512 7X237= 216=7X 
 tpg|BK006948.2| 196420 + tpg|BK006948.2| 196560 - INS GATCCCTACAGGGCTGATACTGGGAAAGATGGTCAAATGGGGACCGTTGCGACCGTTCCTTTCCCAAGAAACAATTGATAATTGGAGTGTTCTCTACAAACACGTACGTTATGGGAATATTCAAGGCGTGAGTCTCTGGCTGAGACAAAACGAGCGTCATTTGTGTGCAAGACAGTTACTGATCGT tpg|BK006948.2|:196034-196946 7X6=87S 89S4=7X 
 tpg|BK006948.2| 198295 + tpg|BK006948.2| 198888 - INS ATAGTAAGATTCCGATTTTTGTTCACTAACTGTGGAAATCTGAGATGAGTTCTTATAGTGGCCACCAGGTTGGACCGGCGTTGGTAATATTTCTTCGGTTAAAAGATCCCCCTCGCCATCACCTTCTTCGATGAACAACCTTGACCTAGGACGGTCCTTACTTCTGGGCGGAATAGTTGGAT tpg|BK006948.2|:197917-199266 7X6=85S 85S6=7X 
 tpg|BK006939.2| 259175 + tpg|BK006939.2| 259903 - INS GCTGTAATGCGTATCTAAGGTAAAACACGTTGAATTAAAAAAGATCTCCTTATTTCGCTAATACCCCTGAAGTCCAACTTTTGGTTAGCCGAGATCTTAGCCGAATGAGATTGTGAAATGCAACCCAAAGTGACCGTTGTTGCTAGCTAGCATATGAATGAATCTAAGAACTGGAAAGGCAAGTTAAGGGCCAAAAATAATGACTTGAATATTTTGCAGTATCTACGTTGAATTAAAGTATTCTTCGTAAGCGGTACTTTTCACTTGCTACTTGTCACCTTATTACCTATGTGCTGAGAGGGTAATGGTACGATGTTCCTTTTTGACAC tpg|BK006939.2|:258503-260575 7X255= 10S294=7X 
 tpg|BK006948.2| 129935 + tpg|BK006948.2| 130220 - INS TTTTGGTATAAAATCAACGCCAAATCCATGCAGGCAATGCCAAGCGGAAGCGATAGAAAACTGGTGAAGAAATCAGTCAACACACTTGGCAAATCGCATCTAGTGACTCAAAGGTCAGCTTCAAGTCCCTCTGTTGAGGAAACTACTCATTCAACCCTATACAATAACAATACTCACGCTTCTACTGAAAGTGAAATATCAATAAAGAAGAGACCCACTGATGAAAGAACAGCGCAGATA tpg|BK006948.2|:129441-130714 13S89=25S 113S7=7X 
 tpg|BK006948.2| 757967 + tpg|BK006948.2| 757621 - INS GAAATAGATATTGTACGTTATTGAATAGTTCTAATATGCAGCAAGTTACTGGTAAGCTTTGTTTTACCCTTGAGTTCGATACTCAGTTTACTTCCTCCATCGGAGGTTGAAATGCGCCTTGTCATACGGCCAAAAAATGCCATGTAAGAAGATGACACTTTCTGCATTTTGAGTATATTTAAGGGCCTATAATTTTCTTCCAACTTTCTCAAGACAAGCATATTGTGTACTTTCGGTTTAGCAAGCCTTTTTACTTCGTTAACACAAGGCGATGCTAACGTGTGTTTACTGTTTTAGAAGATCGGCATTTATCAAATGTAAGGACAATGAGACATGGTTGACCAATTAGTTCTTCTCAGATAGGAGTTCTAGTTCTTCTGCATACTACTTAGTCCTCTTCTGTCGTTGACATTCAATTGCTTGTGCATTTCTAACATGAAATAGTGGTACTACGAATGCTATTATTCTATGCCAGGCAAATTCCTCTGGAACTTTTTTTTTTTCAGTTTTTTCGTGGTGAGCTTTTTTTGCCTGTCTATCTCGAAAGATCTTGTTGTTGATGACTCAGTGCAGTCGCGATC tpg|BK006948.2|:756445-759143 7X6=202S 563=7X 
 tpg|BK006939.2| 394949 + tpg|BK006939.2| 395424 - INS CCTTAATTGTCTACATGGACAACAAAAGACGTGCCCACATAACGTCATGAGGGCTGTCTCTGGAGGTTCAAAACAAATCGGGCAGCGATAGTCCTTGGCTGCACCATACTCTTTGGGTGCTTCTTTGGTTTCCTCCTGAAAGTCGTCATCTGATATTTGCAACACTTGTTGCTCTTCAGCGTCTAAGTCTATGGCATCTGCAGTTAAATCAACAGTTTGTTCCTTACTATTTGTTCCAGGTTTCGTTGTCGGCGGTGCTGCGTCAAGCATCGGGGAAGCACTCGGAGTGTTTGCTGTTTGTGAAAGAACGTCCATTGTGTGCAATTCTTCAACATTATTCGGTAATGTGATATTGTTACCAGAACTTGCTTCTGGCTCTTCGGTATGCATTGTTTCCCTGTCATGATTCCCAGAATCGTTGTTACTGGTGTTATGGTCGCTACCTGGATCTTCTTCAAGTGCTCTAAAGAGAGATAAATCATCATC tpg|BK006939.2|:393963-396410 7X191= 326=1X144=7X 
 tpg|BK006948.2| 1041714 + tpg|BK006948.2| 1041754 - INS CGACCTTTTGGACGTGGGTCCATGGACGAGCACCAGCAATGTATTGCACTTTGTTTTCGGAGAAAGTAGAGTATTCGTTGACGATTTGTTCCAAGGACTTGAAGTTGACCTTAGCACTGGAAATATCAGCGACTTGTTCGGAGGTGATACCAGTTTCAGAGATGATACAACCCTTGGAGTCAGATAGGGAAACGACAGTACCACCTAGCTCAATAACCTTCAAGGCAGCGTATTGAGCAACGTTACCACTACC tpg|BK006948.2|:1041194-1042274 7X154=35S 1S1=319S 
 tpg|BK006948.2| 1040071 + tpg|BK006948.2| 1040457 - INS ACACATTTACCAGTCCGCAGCCGCAGGCTTGAAAAAAGTGACTTTGGAGCTGGGTGGTAAATCACCAAACATTGTCTTCGCGGACGCCGAGTTGAAAAAAGCCGTGCAAAACATTATCCTTGGTATCTACTACAATTCTGGTGAGGTCTGTTG tpg|BK006948.2|:1039751-1040777 7X117=15S 3S1=186S 
 tpg|BK006939.2| 560896 + tpg|BK006939.2| 560477 - INS TTCTTGTATGTGTCTCTGGATAAAAGTATGTCACTGAATTGAAGACTACTGAACCATGGCAGCTAATACAATCACGCCCATCCAGAAAAGTGTCGTGTGGCGAAAATTCTTGTTCACGTTGAACAGAGGGTACTGATTTCAAAGTGCTCTTAAGTCGTAATGACGGCCCTAATAATGATTTCCAGACCCTTTGGAAGGAGTTTCTTCTTTAAGTACTGCCCTCCCTGATCTATATTTGTAGGAAATTTTTAAAGTACCTAGCCTTTTTCTCAGTCACGGCTGTAGAGTGTACACAG tpg|BK006939.2|:559871-561502 7X199= 4S86=1X187=7X 
 tpg|BK006948.2| 413745 + tpg|BK006948.2| 414330 - INS GAAATGGCAACACCTTTTCTGCCGAATCTACCGGTTCTACCGATTCTGTGAATGTAAGTAGCTGGATCTGCTTGTCCGTTAGCAAGCGTTGGAAGATCATAGTTGACAACCATTGAGACAGTAGGAATATCAATACCACGGGCCAGGACATTAGTAGTAATCAAAACTTTGGATCTACCCTCTCTGAAGTCGTCTATTAATCTGTCTCTTTCTTGTGTCTGTAAATCAC tpg|BK006948.2|:413273-414802 7X208=6S 6S1=369S 
 tpg|BK006948.2| 756496 + tpg|BK006948.2| 756704 - INS GGATGTTGTATCAATTTCCACACATTGCTTTAAGCATGATGAATATAGTAAGATATATTACCATCTAAGTTAGCTATTATTGGATGGTTCAACTCCATCAACGTGTGAGTTCCGTTTTTCTTTAATATATCCCAAATGTAGTCATAGAGTGGTTCCTGAACGGGCCTCAACACAGTGCTATTATGGAAGGGGATGTTGTATGGGTTAGTTAATTCTGTAATTCTTAAACGCGGGAACCTTAAGTTCAATTCTGTTCTTAAGGAC tpg|BK006948.2|:755954-757246 7X6=195S 9S231=7X 
 tpg|BK006939.2| 274592 + tpg|BK006939.2| 275229 - INS CTGCCTATCCCTCATCTCTGTCCACTATCGCTAATAATGTTCCCAACATGTATACTATTGCTTTATCGGTGCAAGCCACGTGGGAACCTCTTGCGAAAGTCCCAAGAGTTATTTGGACTTTATTAGGCAATGCGGCCGCACTGGGTATTGCCATTCCTGCCTGCTACTATTTTTCTACCTTCATGAATTACTTCATGGATTCCATAGGTTATTATTTGGCTATTTATAT tpg|BK006939.2|:274120-275701 21S52=48S 108S7=7X 
 tpg|BK006939.2| 194013 + tpg|BK006939.2| 194345 - INS AAGATATACCATATATTACGATCCCTGCGCCCGGCGTGCTCCACATTAAGTAAATGTCTGGAGTAAAATGAAGTCCGCCAATTCAGTCACAAAACATGACTACTGCCTCGTTCGCGATTTCTTCTTCCCTTACTTCATCATGTTCAAGCCCCCTCAGCTGCGCCCAAATGATTCTTCTTATCCTCTTGCATACTGCACCGAAAAAAAAAGTTAATAAGCAGCAGGATTTATAGGCGCGTGCGTGCAGCCTTAGACTGAAGGGGTGGAAAAACTTTAGGTAGGTTTGGTTCTCACTACCCAAAGAGCAATCGATAGGTATAAAAG tpg|BK006939.2|:193351-195007 7X232=51S 2S1=223S 
 tpg|BK006939.2| 13240 + tpg|BK006939.2| 13625 - INS TTACGCCTTGAGAAAACGTAAGGTTCTACATAAATTATTGAGAAAGACTTATTTGAAGATATCGAGAGTCTATCATGCCCTTTGCACAACAAAACTAATGTCAGCTTGCCCTTGCAACATCGTTATACTCCCAGTCGAGATTTTGAAGAATTCATCTAAAGATACTAAGTATAGCTTGTATACAACAATTAATCGAGGATATGATGTCCCAAGACTCAAATATGGCATCATAGTTAGCCCTCGAGTGCACAGCCTTGAGACTTTATTCAGTGATCTGGGCTTTGACAAGAATATAGAGAAATCCTCGCTTTACTTATTATTAAATGATCCTACCTTAGCATACCCTAATTTCCATGAACATTTTGAACAGCTTAAAGGTGAAACAAACAAAGATTTATCTCTACCGACATATTAT tpg|BK006939.2|:12396-14469 7X334= 403=7X 
 tpg|BK006948.2| 95220 + tpg|BK006948.2| 95930 - INS GTTTAGTTCAGCGCCTCTGGGGTGTTTAAAACTCTTGAGGTGACGTTCGTTAACTTATTAACGTCAAGATCTACTTGATCGCTGTTCTTTTTCAAAATCGCGTCCGCTGCATTGAAGTTTGGATTATATCCTGAACTTGGGCCCTCCCTTGTCTCCAGCTCCACATCGTGATCTCTCGTAGATTGCGCTTCGTGATCCTTTGAGAACAGGAACCTCTTGGAG tpg|BK006948.2|:94762-96388 7X5=185S 209=7X 
 tpg|BK006948.2| 259633 + tpg|BK006948.2| 260196 - INS TATATATGGTGGTAAACACGCATATACTGTATGCCATGTATTTACCATTACATAGTTATTTACGCACTCTATAAAAAGTTAACATTGCATTTTAATAAATTCCTTAAATTACTCTAATTAGGATGGTAGCCCTACCTTTTTTTTTTTTGGCACACATGGTCAACTTTT tpg|BK006948.2|:259283-260546 7X6=78S 79S5=7X 
 tpg|BK006939.2| 16775 + tpg|BK006939.2| 17506 - INS ATATTGTCCACAGTCATCTAAAAGAATGACCATTTCGACGACTTAGTTCGGAAAATATTTCCAGCGGATGACACCACTTGCCACAGTTGGTGACCGCCAAATCTAAGTCACACGCGGAAACTGAAAGGTTGTGAGTATATAA tpg|BK006939.2|:16477-17804 7X6=65S 67S4=7X 
 tpg|BK006939.2| 485594 + tpg|BK006939.2| 486166 - INS TATACCTAAAAAATTTGTTGATGTTACGTGATTCCATACAGAACTTTAATATTCAATATACAGTTAATGAAACTTATCTGGATTTTTCTGGTGTTGAGGGGTTTTTCAAATCACTTAAAGAAAATGGTAGAAACGTTTTGAAAAAGACAAAGTCATCTTCAATATTGACCCTGGCAAGAG tpg|BK006939.2|:485220-486540 7X6=84S 84S6=7X 
 tpg|BK006939.2| 301650 + tpg|BK006939.2| 301894 - INS TGGTTGATTTAGGTATTTGGGATGAGGGTATGAAACAGTATCTGATTACACAAAATGGCTCCATTCAAGGCTTACCAAACGTTCCACAAGAATTGAAGGACTTATACAAGACTGTTTGGGAAATTTCACAAAAGACTATCATTAACATGGCAGCCGATCGTTCTGTCTATATTGATCAATCTCATTCTTTGAATTTGTTCTTACGTGCCCCAACTATGGGTAAACTAACAAGTATGCATTTTTACGGATGGAAGAAGGGATTGAAGACCGGTATGTACTATTTGAGAACCCAAGCTGCATCTGCTGCAATTCAATTTACTATTGATCAGAAGATTGCGGATCAAGCTACAGAAAACGTTGCTGATATTTCCA tpg|BK006939.2|:300892-302652 7X3=293S 186=7X 
 tpg|BK006948.2| 803688 + tpg|BK006948.2| 803817 - INS TACGTCAAACAGGCCACCAAGCAATAGACAAGTGCTACTGCAACAAAGGAGGGATCAAGAGTTAAAAGAATTTAAGGCGGGGTTTCTCTGTCCAGACTTGAGTGATGCGAAGAATATGGAATTTCTAAGAAACTGGAATGGCACTTTTGGCCTTTTGAATACTCTAAGATTGATCAGAATTAATGATAAAGGTGAACAAGTCGTTGGAGGAAATGAATAAGAAGTGTCGCAGAGGAATCTTTATGGTTTATATGC tpg|BK006948.2|:803164-804341 7X195=1X9=1X17= 128=7X 
 tpg|BK006939.2| 231182 + tpg|BK006939.2| 231185 - INS AACGCATCCTCACCAAGAATTATATCGTCCGCAAACTTTAACGCAAATAGTCCTCTACAGCAGAATCTATTATCAAATTCTTTCCAACGTCAAGGAATGAATATACCAAGAAGAAAGATGTCGCGCAATGCATCGTACTCCTCATCGTTTATGGCTGCGTCTTTGCAACAACTGCACGAACAGCAACAAGTGGACGTGAATTCCAACACAAACACGAATTCGAATAGACAGAATTGGAATTCAAGCAATAGCGTTTCAACAAATTCAAGATCATCAAATTTTGTCTCTCAAAAGCCAAATTTTGATATTTTTAATACTCCTGTAGATTCACCGAGTGTCTCAAGACCTTCTTCAAGAAAATCACATACCTCATTGTTATCAC tpg|BK006939.2|:230404-231963 7X203= 191=7X 
 tpg|BK006948.2| 546890 + tpg|BK006948.2| 547000 - INS GTTTAATGGTGCCCAGTTAAAGGCGGTAACTGTGGAGGCAGGTATGATTGCCTTAAGGAATGGGCAATCTTCCGTTAAACACGAAGATTTCGTTGAGGGTATAAGTGAAGTTCAAGCAAGAAAATCGAAATCGGTATCCTTTTATGCATAAAAATAATAATATTTTGATTTATCA tpg|BK006948.2|:546526-547364 7X5=82S 81S7=7X 
 tpg|BK006939.2| 84508 + tpg|BK006939.2| 83902 - INS CCAAACCAGATGAGCCCTGGCCATCAGCTTTCTTCTGGGGCCCTGGGCGCCAAACCCGTGACGATCAGAAAAGGACTGACCAATGATTTGGCCGAAGTCCTTCTCATAGATTTCGATGTTACCAAACCTTTTGGACTTGTCTTGTTGCGATTGCGCCATCTGTAGATTGGATAGTAACACGCCCATGGTGTTATCCGAAGAGTCACTCACCAAAAACGACAGATCAATCAGGTTGTGCGGATATGTCATGGTATTCAGATGGTTAAAAAACATGGGAAGATGCTCAGAAGCATCTCTCAGTGGCACGCAAAACAAGATGCGGTCACCCTGTTGCCAACCATCTTTGTTGCCTTGGTAATTTCGTAGG tpg|BK006939.2|:83154-85256 7X5=291S 356=7X 
 tpg|BK006939.2| 382516 + tpg|BK006939.2| 382955 - INS CCATTATTCTTTTCAACTTGATTCTCATTATCCTTTGCCTTTTCTTTTTCATCTGATATTGACTGTGATCTTCTTCTGTATAAAATGGGAGAGTTTTCAAGAATTTTGGACGGCGTAGACTTTATATCTTTAATGACAGACGACGTCACGAAAGAATTAATATTCGACAAGTCTTCCATAATAGTGTTCATATTTGTAGAATTTGGCTGGTTGGAATGCAGGTATTGACTTTCGTTGACTTCAGAATCTGTTTTAGCTATATTGACATCTGCAGTAGAATCTTC tpg|BK006939.2|:381934-383537 7X2=1I2=1X162=45S 2S1=194S 
 tpg|BK006939.2| 170693 + tpg|BK006939.2| 170647 - INS TCTTGGTCCTCTCCTGATAAGTTAGATGTATTCAAACCTGCTATCTCGTCACTCAAACTGATCGAGTCATTCAAATCGCTTCCACCGAGTGACTCAACTTTGGCAATATTTAGTGGTTTTTTTAATTGGTCATGAGCTCTAGCTGTACTTCTCTCGGGCACGTAAGTACCATTTTGCATAGTAGGGGTGGTTTCTGTTTCTTCCGCCAAAACTGCGTTTAAGTCCTCCAAAAGGTTA tpg|BK006939.2|:170159-171181 7X3=442S 119=7X 
 tpg|BK006948.2| 90577 + tpg|BK006948.2| 90379 - INS TGGCACCTAATTGATGACGCACCAGGTTTATATGTAAACATAATCAAAAACACATCCACAACAGTAATGGCCACGCCCGCTGGAAGGGGCACTTTGATCAGGATATTCAAGGCAATCGCTGTACCAATCACTTCAGCTATATCGGTGGCTATAACGGCACATTCTGCAAAAAAATACAATGTCCAGTTGAGCCACCGTGGTAAATACTCTCTGCAAGCT tpg|BK006948.2|:89927-91029 7X176= 110=7X 
 tpg|BK006939.2| 202695 + tpg|BK006939.2| 202759 - INS CTGCGGCCAGGTTGAAAATTTTGATTTGAACAAACCTTACACAGCATCTGATTTAGAAGACCCTGATTATTCAAGCGATGAGGACGATAACGACGAACCCACCCAAAAAGACTTTGATGACCGTAAAAGAAAACACGAAGAAGACATATTCACTGGCAATGGTATAACTATAAAAAGACATCCGGATAGCAAACACATCTTGATCATCTCCAGGGGCCAATACTATAC tpg|BK006939.2|:202225-203229 172S48= 214=7X 
 tpg|BK006948.2| 853133 + tpg|BK006948.2| 853359 - INS ATAGGAGATTTTCTCCGATCCAGAAAAGGGAATTGGTGGACCTGAAATGCAGTTGCAACATCTTAGGCAACTTCAAAACTATTTTTCGAGGTGGTGGTAATCCAAATGGGGACATTTTCGATTGGGAACTCGGAAAGCACGGTATTGAACTGTATTTTAAGCATCCCAAAACAGGCACCACATGTAGCGCAACCTTTTTACCTGATGTTATGCCTGAGCAACATTGGAATAAAG tpg|BK006948.2|:852651-853841 7X130=45S 1S1=160S 
 tpg|BK006939.2| 182546 + tpg|BK006939.2| 183131 - INS ATAATGCTTTGAACGAATTTAAAAACGTCAAAATAGTTACTGGGAACCCGGTTACGCAAATAATGAAACGCCCTGCTAACGAAACGACAATCGGATTGAAAGCGAAATCTGGCGACCAATACGAAACATTTGACCATTTAAGACTTACGATAACACCTCCCAAAATCGCTAAATTGCTACCGAAGGATCAAAATTCATTATCCAAGTTATTAGATGAGATACAATCAAACACAATAATTTTAGTTAATTATTATTTGCCAAACAAAGA tpg|BK006939.2|:181996-183681 7X1=1I233=14S 1S1=192S 
 tpg|BK006948.2| 560312 + tpg|BK006948.2| 559857 - INS GCCATGACAATATTTCTATTGTTTTTTTTCCTGAAAATCCCGTATATGAAAAATTATACAGTTGCTTAAAAGTTAGGGAAATATAGACAGAGTACGTACAAAGGATTACTGCATTCAAGACATTATGTTAGATCCATCATCTAGCACATCTCTCCAATCTTTCAGTTTGTACTGCATGTTTTTGGGATGATATTGGGGGTAGAATGTCTCAATGACCTTCAATAATTCGTCATGAAAAATTT tpg|BK006948.2|:559359-560810 7X5=106S 227=7X 
 tpg|BK006948.2| 565292 + tpg|BK006948.2| 565953 - INS AAATAGCATATGCTGACATCCTATGTGGAGTTCTATGAGCAGAGACTATTGTCACTTCAAATGGAACGCCAAAATCTTTTAAAACCGCACATGCGGCAGACATTACCGGCAAGTCAGAGTCTGATCCCATGATGATTCCAACCAATGGTTTGACCATTGCTTCCAAGTCCAACTTTTGAGCGACAGAGATTTTGATTGGAATATCAGTTCTACCTGTAA tpg|BK006948.2|:564840-566405 7X2=406S 110=7X 
 tpg|BK006948.2| 602706 + tpg|BK006948.2| 603009 - INS TCAAATCAGCCTCAGTATCAACGCACCAAAACTGCAAGTGCATCAAGCACTTCCTAATATCCGCATTATTTTGTTTTACAACATCGCGAAGCCAGTCGTCACAAACTTCGATTTCAAGGGACTTTAAATATTTTGTTAGAAACGCATAGACTGTGGATGTACTAATTTTCTTAGTATGAAACAAAGAGTTTTGTTCACTTGCCAAGGCAATAAGTTCACTAGGAACTAGTGACAAATCCTTACAAG tpg|BK006948.2|:602200-603515 7X6=117S 118S5=7X 
 tpg|BK006948.2| 246009 + tpg|BK006948.2| 246123 - INS GGTTGATGATCCTAAACTGGTGTTTAAACAGGTAGTCGCTAGTATAAAGCATTTACATGACCAAGGAATTGTTCATAGAGACATAAAGGACGAAAATGTTATTGTTGATTCTCATGGCTTTGTAAAATTAATCGATTTCGGTTCGGCTGCCTATATCAAGAGTGGACCATTCGATGTTTTTGTGGGAACAATGGACTATGCTGCACCTGAAGTCCTTGGTGGTTCCTCTTACAAAGGTAAACCA tpg|BK006948.2|:245507-246625 7X206= 229=7X 
 tpg|BK006948.2| 313421 + tpg|BK006948.2| 314150 - INS CCTCAGGGTTCACTCTTTCCAAACGAATCTGTTTCTTTTCTTGGGAAGTCAGTTGCTTTTTCTGTTCTTTTTGTAACTGGAAGTAATCAAACATTTTGGTGAAATCGCAACGAGAAAATTCCTTTATCTCAATTCCATTGAGGGGACCACCACTTTCTTTCAGTACTTGCAAGAAATCATTGAAGAAGTTCTTTTGGAAAACAGGATTTTTGGCATGATCACTCTCTAATAGGGCAGCAAAGAACCCGGCTACTTCTTCAGCTTGCGGAGGTAAATCTACTGGCTTCCCATCGTAATATAATTTGATGTGAGATGGTAAGGGCTGGTATGGTGGAGGG tpg|BK006948.2|:312731-314840 19S157= 86=90S 
 tpg|BK006939.2| 478032 + tpg|BK006939.2| 478169 - INS ATTTGACACTACTGATGATCTATTTGTGGAAAAGGAGGCCCTTGAATCTCTTCTATTCCTTGCTGAATTATTGCTTTCCATAACACTACCTAGAGAAGGCGTTTGACCGGTGTTCTTATTGATATTATAGCTATGATCGTTGTCACTATGAGTACCTGAGATAATAACAGACTTCCTATTCTTTTTCGGAACGGCCTGAT tpg|BK006939.2|:477618-478583 7X5=95S 95S5=7X 
 tpg|BK006939.2| 189687 + tpg|BK006939.2| 189867 - INS AATCATGTCTGTGTAACCTTTTTGAAATCATCATGAGCACCGCTAGTCACCGATGGAAAATGTAGCTCCTCAGAAACACGGCCACCAAGAGCCATGATCATTCTATGTCTGAATTGCTCCTCAGATATCAAATATTGATCCGGTGGTAGGTACTGGGCATAGCCTAAAGCACCTTGTCCACGCGGGATGATGC tpg|BK006939.2|:189287-190267 241S32= 97=7X 
 tpg|BK006939.2| 431478 + tpg|BK006939.2| 431967 - INS ATCTATAGTACTAAAGCTTTTGCGGTTGTTATTCAATTGAGGTAGATACCTGGCAAAACATTTCTTGTGAGCACAACCTCAATTAAAGTTAGACAAGTAGGTGCACTATTGGTTGCTTGTTGGCTCATCTCGTTGAGGAATGTAATAACTACTTGTTATTAACCTGTTTTTGTGCCATCTATAGTGGAGAGCTTATTGCAATTTGTTTTTTATTTCTTGACTGCATATATC tpg|BK006939.2|:431002-432443 7X205= 116=7X 
 tpg|BK006948.2| 197328 + tpg|BK006948.2| 197395 - INS GGGCATACTCGTTGTCTTCCCTTTGTCACACTCAACAGTTGATTTAGTGTGTCGATATCAAAGGATCGCAATTCCTTCACAGATTTTTTTTTATTGAGCTTTTTTTTCGTATCCTTCTTGAGTTTAGTTTTCTTGGGCGTTTCCTCAATGATGTCCTCGTACATGTCATCATCTTGTTTGTTTGTCGAAGTAGAGGTATGATTTGCCCTATCATGAATAGCCTTCAATGTGTCGTCACGTTTCAAATTCGATGTAACTCTGCTATCCTCATTGGGTGTGCTGGGCAATGGTCTTGTCAAGTAAGTCTCTTCCTCTGGAGGCATACTCGTTGCCGCAGAATAGTAAGATTCCGATTTTTGTTCACTAACTGTGGAAATCTGAGATGAGTTCTTATAGTGGCCACCAGGTTGGACCGGCGTTGGTAATATTTCTTCGGTTAAAAGATCCCCCTCGCCATCACCTTCTTCGATGAACAACCTTGACCTAGGACGGTCCTTACTTCTGGGCGGAATAGTTGGATTGTAGTCATTGGTTTCAGAACGTATTGGGTTTATCGCTTTGGGTGCTTCGTTGGTGGTTGTATACAACTCGGGTATGACACTGGAAACAATTGAAAGC tpg|BK006948.2|:196078-198645 7X4=155S 599=7X 
 tpg|BK006948.2| 454554 + tpg|BK006948.2| 455193 - INS ATTCAATTGAATCAATTGGTCAAATATCTACAAATGAAGAAAGAAAAGACAATGAGCTTTTAGAGACCACAGCTTCATTTGCGGACAAGATAGACTTGGATAGTGCGCCAGAATGGAAAGACCCTGGTTTGTCGGTGGCTGGTAATCCGCAACTAGAGGAGCATGACAATTCCAAAGCTGACGAT tpg|BK006948.2|:454170-455577 7X5=87S 86S7=7X 
 tpg|BK006939.2| 371583 + tpg|BK006939.2| 371004 - INS TGGAGTTGAATACCTGCATCCCCTTCTAGTACTTTTTGTATCAACTTTCCTCCGGGTATGCTAGGTATTAGTTTTGTAGGTAGTAAATTTGCTAAGTTTGACTTTGTCAAACATATTTTGTTACTCTTGCTATTGAATAGGTTCTCCGAGCAGTTATATTGTAATTCCCACACGTTGACACCATCAGT tpg|BK006939.2|:370614-371973 7X5=213S 177=7X 
 tpg|BK006948.2| 925260 + tpg|BK006948.2| 925288 - INS CAAATCGGGTGATAACGTATGTAGGGCTAAAATAGATATTGAGTAGGTTACAATTAATTATTGGCAATTGCACCTAGTGACACATTTACGAAAACGTAGGGCAAAAACTATTACCCGACCCAGGGCTATTTTGTGATTTTTTCCTTTTTTTTGTTTATGATCGCGCTTCTCGAAAAGCCAAATATCAGAAATCCCAAACACGCCTTCATTTGATACGATTCGTAGCCTGCGTTTCAGAGATCTATCAACTT tpg|BK006948.2|:924744-925804 84S82= 236=7X 
 tpg|BK006939.2| 90464 + tpg|BK006939.2| 90704 - INS ATTTCAAAGATTAACTGCCTTGAAGGAATTTAGAACTATGGGTATCAAACCTTATACCATTAACGTGTTTAGAAACAAAAAATGGGTAGCATTGCAAACCAATGAATTGTTACCTATGGATTTAGTGTCTATAACAAGAACCGCCGAGGAGAGCGCAATTCCTTTCGATTTGATCTTGCTCGATTGCTCCGCTA tpg|BK006939.2|:90062-91106 7X142=27S 7S1=119S 
 tpg|BK006939.2| 399249 + tpg|BK006939.2| 399617 - INS CTTCAATTACCTCATTGAGGTCAAGGCTACTGTCGCGAATCAACGGAGAACTTTCGGTAGCAACAGTGGGTTCATCCGCCGATGTAGCACTTATACTTACATTTTCCTCGGCGAAGTGTTGCAAAATCTGATGGATTGAAGCTCTTGCAGGATGACACTGTAGTGGGAACGCCAGCATCACCAACAACACAAT tpg|BK006939.2|:398849-400017 7X96= 182S3=7X 
 tpg|BK006948.2| 874115 + tpg|BK006948.2| 874462 - INS ATATTATATATACATAATAAAAAAGGCACTTTAGACAGAATGAGAATACTAGCAATCACGAATTCCTACTTTTCCTTTCTGTATCCCTAGGCGTTTCACTCGACAAGAATTGATCGTCTTGTACCAATCCAAGCAGATCGATATATACATATATATCTGGATTTCGAGAAGAAGGATATATTATATTGCTTATTTGTCTTTTTATAAAATCTCTCCTAAGTTAAGT tpg|BK006948.2|:873649-874928 182S157= 168=1X43=7X 
 tpg|BK006948.2| 100347 + tpg|BK006948.2| 100793 - INS TTGTATATGATTCTAAAATAATGTGTGAAAAAAAAAATAAAATAAAAAAAAGAGGAAAATAATATAGAATAACTATTAAGTTTCATTAAAAAAAAACCATTTGAATATACGACCAAAAACGTTACGCTTTCATAAAGTGTGAATAAGCAAGGGAACTATACTTGAAATATGGGGGCAAAGAGTGTAACAG tpg|BK006948.2|:99953-101187 7X7=88S 89S6=7X 
 tpg|BK006948.2| 1001324 + tpg|BK006948.2| 1001626 - INS CCAGGAGAAATGCTTCCTTCACGATGGGATCTTTCTTGAACTTTTTAGGAAGTTCTTCTTCCCAAAATTCCTTTAAATGGTTGAAATTTCCAGAATCAGTTAGTGCGTTAACTAGCGTCGCATAAGATGTGTTTTTAATATTATCTCCTGGTTTGATAACACTGTTCCAGACTGCTAGAATGC tpg|BK006948.2|:1000944-1002006 7X24=67S 8S1=274S 
 tpg|BK006948.2| 922270 + tpg|BK006948.2| 921898 - INS CTTTGTGTGTAGTCACTCCGCCTTCCAAAGTTAAGTTTTCCAGAACTTCCCACCACTTAGAGAATTTTGGGTTAATCAACAACGTTTCCATAGCGTTGCAACCAGCTGGGTAGTTAGTCTTTGCATCCAAACTAATTCTGTTTGCCTTAATCAAATCTGCGTCTTCATCCAAGTAAATTGAGCAGATACCATCCGCATGACCCAACACGGGAATTTTTGTAGTGTCCTTGATTTTTCTGACTAAGGCATTGGAACCACGAGGAACAACTAAGTCGATGTACTCATCTTGATCCAACAAGTCGGAAACATCCTGTCTGGTTTCGATCAATTGCAC tpg|BK006948.2|:921216-922952 7X152= 119=1X194=7X 
 tpg|BK006939.2| 251824 + tpg|BK006939.2| 252113 - INS CAACCAAAGGTTACATACCTGGTGAAGAAGAAGCGTGGGTCCGTAACAACACATCCACTTTGGCGCAGATTGAATCTAATGTCCTAGAAGATTTTGAATTTCCAAAGGACGAGAGAAATATTTTATCATTTCATGAAGTGAAGCACTTTGAAAAAATGCTCAAGGGCGATGCTGGCGCAAAAACTGATAACACACCTAAAGAATCTATGACTAGTGTGATTTCTGATTCGGTTAAGTTGTCTGAAGCCGAGTTCACCTATCTATCTCAATACATCTCTCCTGAACATTTAAGCTCGAAAGG tpg|BK006939.2|:251208-252729 13S245=21S 24S5=7X 
 tpg|BK006948.2| 274977 + tpg|BK006948.2| 274671 - INS ATGATCAGCTCCCCGATTTAGTTCTTTCTATGATCAGCGACCCTGCAGCTGCTCAGTTGGGATGGGTAATAAGCTTGATATGCGACCCTTTATTAAACCAAAGCATGATACATGCAAATCGTTCTTTTGTTCTGATTGAGACACTAAGAAATGTGTTACAAAAAATTGAAAACTCCCCTCATTTAGATTACCACCAACCAGTAAACAGTTCATTAGAGTTTATCTCCAAATTTATTGTTGAAATGAAAAGGCATATGTGTGATG tpg|BK006948.2|:274129-275519 7X293= 132=7X 
 tpg|BK006939.2| 469574 + tpg|BK006939.2| 470117 - INS TCCGCTCACTTCATGCCAACCATTTTCTTCGGTAGAGTCATCATTGATCACGCCATATTTTTCTATCAACTCCTTCAGTCTAGGACTAGCATTTTTGATAAACTCTGCTTTTCCATAACGTGACAAATTTCTAATAAAGAAAACTTTCAATTGTTCATCATTAATACTTTGCAGCATATTTTGAATTTCATTATCGGTTAAGCCATCAATTGCAGAAATTAATTC tpg|BK006939.2|:469110-470581 7X179=17S 2S1=269S 
 tpg|BK006939.2| 221706 + tpg|BK006939.2| 221770 - INS GTGTAGATGGTAGAAAGTCTAAGGAGTCATCACTTGACCTTTGAGAACTATTATTAGTATTGCCACTGAAGTTGCTATGTCGCTTGGGGCTTTCATCAAACGACGTGGACTTCTTATGGGCTTTTATGAAAGACCGCATGATGAAATATTCCAGTT tpg|BK006939.2|:221380-222096 7X5=73S 74S4=7X 
 tpg|BK006948.2| 837532 + tpg|BK006948.2| 837546 - INS ACTATACGTTTTGAAACTGAATGCATGAACGCTATTGAAGATATTCACCGGAGGGGTAAGATACCCATCGTTGTTGGGGGTACTCATTATTATTTGCAGACTCTTTTCAATAAGCGGGTCGATACGAAATCATCCGAACGTAAGCTCACAAGGAAGCAGCTCGATATTTTGGAATCGACTGACCCTGATG tpg|BK006948.2|:837138-837940 7X9=86S 91S4=7X 
 tpg|BK006948.2| 111155 + tpg|BK006948.2| 111776 - INS GAATATTTTGTTTGATACGTAACAAGCTCATACAAACCAAGCCAAGAAAAAGAAGACGACTAATCTATTTATAACAAAGATATTTGTTCACTATAATGCAATATAGTTCGAGGTTCCTAGAAT tpg|BK006948.2|:110895-112036 7X30=31S 4S1=165S 
 tpg|BK006948.2| 786310 + tpg|BK006948.2| 786700 - INS GTCTATACCCTCACTGAAGAACATTGCTTTATTATGCATAAAGGAAAAAAAAATTACCCTAATTTGATTACTTCGTTTCGGATGAATTTGAAAAAAATCATATTGAACCATGACCGATTTAGCCATCCAGAAAGATGGAAAACAAACGCACTCTTAAGGTTCACCTTCGTGTATATAAAATTTCTCTTCGACTTGATGATAATCAAAAATCCATTAAGGATGGTTGGAAAAACTTATCGAGACGCTGTTACTGCGCTAAACTC tpg|BK006948.2|:785770-787240 7X187= 247=7X 
 tpg|BK006939.2| 518959 + tpg|BK006939.2| 519443 - INS GTTATGTCTAGCCCGAAAAAAGTTTTGCTAGAGGATCCCAGAGACAACCATACTAAGGCGAAGAAGAGTAGTAGAAAGAAATCAGGTGAAATGGTCTTCGTCAATTATACTGTACAGGACACGGCTAACGAAAATGATACTGACTTGCAAACCCAGCCGGTTTCTGTGCCAGCACCAAAGGCGAAATTAAAGAAGAAATCCTACAAAAGGAGAATGCTGAAGATATTTGGATCGTCAAAGAACGAACACATAGAGGACATCGTTGAA tpg|BK006939.2|:518411-519991 7X4=155S 69=1X64=7X 
 tpg|BK006939.2| 37147 + tpg|BK006939.2| 37179 - INS TCTCTTCTGTCTTGCCTTCTAATGAATAACTGAGTATTCTTTACATACTTTGTTTTTATTAACCACTAGTTTGAATATATATTCGACTGAAAGGCAATATCAACTATTCAATCTTTAACATTTTTCTCGAGCCCT tpg|BK006939.2|:36863-37463 7X8=59S 65S3=7X 
 tpg|BK006939.2| 260746 + tpg|BK006939.2| 260911 - INS GGGCTAGATTAGCTGATTTAAATCACTGCAAGTAAGGAACATCGCTCTTGTTTCTGTTCATGACTGTTCTATGAGCACCAAAGTAGAAAACGAAAATGAAAGCGAAAATACTCAAAAAAATCTCTAAATCTTGCATTGTAGTGTGTACTGTGTAGTAAAGCTATTGTTTGTTTTTATTATTTCTATGTAGAATTC tpg|BK006939.2|:260342-261315 100S112= 98=7X 
 tpg|BK006939.2| 248333 + tpg|BK006939.2| 247594 - INS GTACCCTCAGTGCTCTCATCTGCTTTTTCGGTTTCAGTGGCTGCTGTACCCTCCTCATCTTCCTTTCCAAACATTTCTGTTGCCTCGTTTAGCTCTTTGAACAAAGAAAAGTCTCCAATCCAATCTTTGAAGCCATCACCACCGAATATTGCTGTAAAGTATTCAGAAGCATCTTCAAATCCTTGCTGAGGAACAGCATCCTCCTTACCAAACTGGTCATACTTGGAACGAAGCCCTGGATCACTTAAGACTTGGTAGGCCTCGCCTACGGCTTGAAAC tpg|BK006939.2|:247022-248905 7X6=391S 140=7X 
 tpg|BK006939.2| 82804 + tpg|BK006939.2| 83060 - INS ACCTTGTGTTTCTATCAGGGTCGAAGTCTAATGGAACTTCTTTAGGATGTTTTTTCTTGTTCTTGTCGTTGTCATCAAGAGGTTTCCCCTGCGGGTTGCCGTCGAGCTGTTGTTGCTGTTGCTGTTGCTGCTGCTGCTGTTGTTGTTGTTGTTGCTGTTGTTGTTGTTGTTGGTTGTTTGGTGAGACAAAGTCACCCTTTGAGTCCACCAGCTCCGAGCCATCTCCCTCTTCAGACCAGTCTACAGT tpg|BK006939.2|:82296-83568 74S208= 124=7X 
 tpg|BK006948.2| 491920 + tpg|BK006948.2| 491888 - INS AAGTGAAAGGACCACCATGTCCATCAAAAATTCCAAAAAAATACAAATCCTTCTCTATGGACTTGCCATCCTCACTTTCTATCGGAATGGTAATGATTTGTTCTACGTGATCGTCTTCTATTGGATGGTTAGAGGGCAACTGTGCCACATCATACCTGAATATACCAGTGCCACGGTTAACAAAATGGCTTTCCTCTCTATCATGTAGTTTAGCCTCTATTTTAGAAT tpg|BK006948.2|:491418-492390 7X162=37S 1=166S 
 tpg|BK006948.2| 339358 + tpg|BK006948.2| 338763 - INS CTTCTTCGACGAATTTACCTGAAAAAAAGAAAAAGTAAACTACAGTCCCTATTTAAGTATTTCGCAAGTCATCTCAAAGTAAAAATAAAATTCCTGGTAACACTCATCCTAGATAGAGCTATATTTGTATCTACATAACATGTATTGCATTAAAGGCTTATTTCAGTCCACTATTGCTTGTTCTCATTGTCTGGTGTTTCATCTGTAGATTGGGCACCTGCTCCACCAAAAAGATTGCCTGCCATGTTTCTGAG tpg|BK006948.2|:338241-339880 7X4=222S 127=7X 
 tpg|BK006939.2| 62260 + tpg|BK006939.2| 62428 - INS TTCTAGTACATAATTATGTAGCACTATCGACTTCCTTTTGGGCATTTCTATAATCTCGAGGAAATCTTCTAGTATATCCTGTATACCTAATATTATTGCCTTCAACACAGACGGAATCCCAACAATTATCTCAAAATTCACCCATTTTTCACTCTCAAATCTGAATCTAAGTAAATAGTGGCAGTGAAATCCGGATCAAAATTCAGTAACTTTTGTGATATCTCACATTGACATACCACGGTCGGAGGTGAAT tpg|BK006939.2|:61740-62948 7X206= 127=7X 
 tpg|BK006948.2| 655868 + tpg|BK006948.2| 655286 - INS CCGGAAAATATTGTGGGGAGTATGGAAAGTTTGGAAAATTTGTGGGTTTGGATTATATTATCAGATTTCAATGTTTCTTTAAATATTGGGAGATGTTTGGCGATTAACTCATCCTATTTTCAAGTCGATGAATGCGAGAATGGTGAGAGGTTGCCTAAAAATACAAACAATTATTCATCGACGGTTTTTTTCGATCAGTCAAATTCCTGCATGGGCAAGCTTAAAAGGTTTTTAAGATTAGCTCGACCAATGCTAGATCAAATTTATGATAGAAGCGCATTTCCAGACTTAGCCGAAAATTGTAAAAAACTAAGAAACTTTGTAGAGACTGAATTCCACCCAATATCATATTACACTGACAGTGAGTTAATATCTAAAGTTCCTTTGTGCGAGATTAAAGTGCTTGCGCAGGTT tpg|BK006948.2|:654444-656710 7X5=335S 207=7X 
 tpg|BK006948.2| 860878 + tpg|BK006948.2| 860849 - INS AATGCCGAGGGCTTCTTTTTCTTCTACAGCCACTACTTCTACGGCGGCCACATTGACTTCCGCGATGGTACTGGATCAGAACAATTCGGAACCGTACGCAGGTGCAACATTCGAAGCCGTGCCAAGTTCTATTGTATCATTCCATCACCCTCATTC tpg|BK006948.2|:860523-861204 7X6=72S 74S4=7X 
 tpg|BK006948.2| 557421 + tpg|BK006948.2| 557883 - INS CCCTCGATTGCAGGCCCTTTTGCATGACCTTCGGGTCTGTAGAATTGAGAAAAATAGTATCGCAAAGTATATCGTCCAAAAGTCTGTCAGAAGTCTTCAGTGGTAGGTTGGTGGCAATATCTGGATACAGTAAGTGTTTTCCATCGTCAACATCTCCAGGGGTAGACTGCTGGTTTATACTTGTCCCGTATAATGGGAGGTCTTCTATAACAGACCCATTTCTGTCAGCATTTTCTTTATCCTGGTTTAGTAGTTGATTATGATGGTTCTCAATTGCTTTTTGAAGTTCATTATCTTCGTTCGGCATTTCCTTATACC tpg|BK006948.2|:556771-558533 7X198=40S 6S1=184S 
 tpg|BK006939.2| 30172 + tpg|BK006939.2| 30552 - INS TTAAAACATCTCTCTTCTTCTGAATACAATTATAATCATACTTATAACGGCCAAGAAAGATGCCTTTGATAGTGCCTCTATGTTTCTCTTCATTGATAACGGAAAGGAAATGAAAGTAGTGACCATTACAATTATGACATTTCGCCTGAGCCAAAAATGTACATTACCATCGTTCTGGCTGAATATAGCTCTGAGTACGTGGGGTATCGTATCCCCAATAATTATGCAATAACCAATACATCCACCAAATGCAAATAACCCGTTTGTAAATAGAATCAGCAATTTCCCTTTTTTACCCATTACATGTTCGACCGTACCC tpg|BK006939.2|:29520-31204 7X202= 5S295=7X 
 tpg|BK006948.2| 590404 + tpg|BK006948.2| 590605 - INS GTACTTTTCATCAGCATCTTGGAAAGTGGTGAAATTTTTCTTCAGCCGTTCAGCAAGAAGCCATCCATGTTTAGAATCGATCTTCCAATCCTGTAGGGGGAAATCACTTTGTAGCAAAAATAGAGCGAAGAGCCTTGTAATATCATCTCCACCATAATCTAACGTAATTGCACTATGTTCCAAAACTGTTCCTTCATCAACACAGGCGATCCTGGTTTCAGCAGCGCCTATATTTACTACGCATGTGGAGGTACTGATCCCGGCACCGTAACAAGTCGCTAATGATTCTTGTATAATAGCGACTGCTTGAAATTGTAACTCGGTGAGTAGAACTCTAATGAACG tpg|BK006948.2|:589702-591307 7X184= 323=7X 
 tpg|BK006939.2| 343765 + tpg|BK006939.2| 344408 - INS GTATTGATGATGCAGATACTGGTTCTGCTGAAACGGAACTCCCACGCTTAATATCTCAAGCAACAGTAGAGAAAGTACCCGAATTGAAGTGGTACAATGATCAGATATCACTGATTACAGAAAAGTTGGAGGACGATGAAGATATTGAGGTTCACGAGGAGCTAATGGATG tpg|BK006939.2|:343409-344764 7X6=79S 82S4=7X 
 tpg|BK006939.2| 108599 + tpg|BK006939.2| 109182 - INS TTTGAATTGAAGTTGGAAAATGGCTTCAATTCCTCTTGTTGAACATTCTGTATCTCTCGCGTATGAATTACCTTCTAAGAATGAGTTCAGGTCCAACAGCAACTCTGTAGTTTCCTCGCTTTTGCTCGATAACAACCTTCCAGGGTTATCAGGAATGAGTGGAGAAGGATTACTAATAGAATGTGCGCCACTTTTTAAAGTGTATTTTATCAAAGGATTTTCCGGGGTTAGAT tpg|BK006939.2|:108119-109662 12S197=12S 14S5=7X 
 tpg|BK006948.2| 661795 + tpg|BK006948.2| 662166 - INS GGGTGGCCCCTCTAAAGTTGAGGAAACATATGATTTTTTGTATCAATTATTTGCCGATAATGACCTAATTCCCATTAGTGCTAAGTATCAGAAGACAATTGCTAAATATATTGCTAAGTTTCGTACCCCCAAGATAGAGAAGCAATATAGGGAAATTGGTGGGGGCTCCCCAATCCGGAAATGGTCTGAGTATCAAGCCACTGAGGTCTGTAA tpg|BK006948.2|:661355-662606 7X69=37S 11S1=26S 
 tpg|BK006948.2| 844178 + tpg|BK006948.2| 844109 - INS GTATTTGGGTGACAGTAACCGCCTACCAGGTTCCCATCTACGGGTTGCGTCCATCGGACCTACCACTAAAAAATATCTGGATGATAATGATGTAACCTCTGATGTGGTCAGTCCAAAACCGGACCCCAAGTCGCTATTAGATGCTATTGAATTATACCAGCGCCATAAATAATATTGATACGTCA tpg|BK006948.2|:843725-844562 7X5=87S 88S5=7X 
 tpg|BK006948.2| 642399 + tpg|BK006948.2| 643070 - INS GGTATACATTAAGCAATTCGAGAACTCTCGAAAAGATTCAGAAGTAGCAAAGCACCCGCCAAGAACCGAATTTCATTTTTATGAATTAGAGATTGAAAATCTCCTTGATAAATTTCCGGAATGTCACAAAAGACATAGAAAGCTATACTCTTATACAGAAGCTAAACAAAACTTGATAGACGCCAAGAGGCCTGAATTGTTGGAGGCCCTTAATAGGTCTGCTATCATTAAAGACGACAAATAGCTAGCACATACATATATATGTATATACG tpg|BK006948.2|:641841-643628 7X195= 136=7X 
 tpg|BK006939.2| 307663 + tpg|BK006939.2| 307737 - INS GGATATGGTACTGAGGAGTATGTTATGTTGATGGAGAACGGTTAAAGTTACATTTCATCAGTTTTTTCCCGTTCTTTTTCACCTTTTGTGAGAAAATTTTACTAACGTTTCGTATATTATTCTTGTAGTACCATTAATTGGAATAAATATACTGGTGATTGTTTATGAATTACTATTGGGATGAACTAAGC tpg|BK006939.2|:307267-308133 7X13=10S 168=3X4S 
 tpg|BK006948.2| 991552 + tpg|BK006948.2| 992041 - INS GTTTATCGCCGCAGGTTCTACAATCACTACTTTCTCATCTGTTAATAAACGCCTTTTTTGACCCCGAATTAATAATCAGATACTCGAGTTTTGCCGCGCTCCAAGAATTATTGGGCAGGTCCAACAAATCTCTTGCGCTAAATCAAAATGACATTGCTTTGATATTG tpg|BK006948.2|:991204-992389 7X5=78S 79S5=7X 
 tpg|BK006948.2| 700810 + tpg|BK006948.2| 701259 - INS GCCGTAGATTGACTATTAGCATCTCTTTTTGAGTATGCTAAGAAGTAGAGGGCTACCTTATTCCCACACACTTTTTACCACGGGCGAAACATTTATTTTCAAGTCCCAGCACAGTGATGGGATGAAGTCCAGGATGCGTCATACGGTCCTATGGCAAACTTCGGGGAAGGTTTAATATGCTGCTTTCAAGCAGGATTAACGGTAATCAACTCCCTAGGCAAATTGGCTCAACTCTGCCTATCTATCCACTGAGGATTTCAAATCCACCGAATGGGAGAATATGTC tpg|BK006948.2|:700226-701843 7X176=37S 2S1=236S 
 tpg|BK006948.2| 465194 + tpg|BK006948.2| 465735 - INS CCAAGAGAAATCGGGAAACTTCACATAAAAGGAAAAGTTTATCCCAAGATTCAATACCCGACGAACCGCAATTGAGAGAAGTCGTCGTCTCAAAGGATTATGGAACTCCAAAAGGGAAAAAAACGGAAGATGAAATACACGAGGATACCGCTCATCTAATGACCACTTC tpg|BK006948.2|:464842-466087 7X92=34S 1=115S 
 tpg|BK006939.2| 217934 + tpg|BK006939.2| 218318 - INS GTCACCTAAGATCATCTCTTTCAGAATCAGAGAAGTTAAAATCCTCTGGAATGCCATTAATTTCATCGATGTCGTAGTGGTCGAAATCAAAAAACTTACTTTTCTGATTGTATTCGTCTTCCTCAGCTTCATCAATGAAAAAGAGATTACTCATTGGTCTGGGGACTTCTGAATCTAAATCGCAATTTAAGTCATGATATTTTAGTGATTGAGACCTAGCTGGCGGCGGAAGAGGGGGGCTATTGAGTACAGC tpg|BK006939.2|:217414-218838 7X164= 127=7X 
 tpg|BK006939.2| 355221 + tpg|BK006939.2| 355944 - INS CATTAACAGAGAAGCTTCACGAAGGCTGTAAAAAAATTATTGTGGGAAGACCGCTTTTAAAGCAAAGCGATTCCTTATCAAAAGCTTCAACTACAGATTGTCAAGCAAATTCGCATTGCCAGTGTGATTCACAAGGCAGTAGGATTACATCAGTGGATGATGATGTCCTTGTTAACCCTGAGAGCTGTAACGATGCTGCCAACAATTCTAATAATAATAAAGAG tpg|BK006939.2|:354759-356406 7X94=18S 1S1=211S 
 tpg|BK006948.2| 929243 + tpg|BK006948.2| 929416 - INS GGATTCGAAGGAGTATGTTTCATTGGTCACAGAACTAAAGGATGATTTCGAAGCTCTAAGTTATAATATATATAACATTTGGCTGAAGAAATTGCAGAAGCAATTGCAAAAAAAGGCCATCAATGCTGTGGTCATCTCCGAATCATTACCAGGTTTCAGCGCGGGAGAAACCAGCGGGTTTTTGAACAAAATTTTTGCTAACACTGAAGAATATACAATGGACGACATTTTGACCTTTTTCAACAGCATATACTGGTGCATGAAATCTTTTCATATTGAGAATGAAGTGTTCCATGCTGTAGTCACAAC tpg|BK006948.2|:928611-930048 9S9=1X86=1X64= 155=7X 
 tpg|BK006948.2| 944986 + tpg|BK006948.2| 944998 - INS CTTAAGCCCTCACAAATCTGTAGGACAA tpg|BK006948.2|:944916-945068 7X4=10S 10S4=7X 
 tpg|BK006939.2| 440965 + tpg|BK006939.2| 441681 - INS TAACAACCCTGTAATGGCTTTCTGGTGGGATGGGATACGTTGAGAATTCTGGCCGAGGAACAAATCCTTCCTCGCGGCTAGACACGGATTGCACGCCCTTTGGGCAAGGGATAGTTCTCTATTCCGCACCGTGCCCTGTTGTGGCAACCGTCTTTCCTCCGTCGTAAATTTGTCCTGGGCAGAGCTGTCTGCCCGGAGGCGGGAGAGTCCGTTCTGAAGTGTCCCGGCTATAATAAATCGATCTTTGCGGGCAGCCCGTTGGCAGGAGGCGTGAGGAATCCGTCTCTCTGTCTGG tpg|BK006939.2|:440361-442285 7X277= 277=7X 
 tpg|BK006939.2| 8134 + tpg|BK006939.2| 8278 - INS AAAAAAATGAACAATAATTAACACGAGAATTTAAACCATACTCGGCCGGATTAGCGATCATTTCGTTAGTAATTAAAATTAACATTTCCATGTGGGACTCTAACTGCTGCATCGCCAAGTTGATAAGCCATGAAATCACCAATATCAAAGATAGCAATCCAACTGGAAAAATTATTCTCGGCATATGGG tpg|BK006939.2|:7742-8670 7X6=88S 91S4=7X 
 tpg|BK006948.2| 85389 + tpg|BK006948.2| 85981 - INS TTTCATATCAATCTTTCCTTCAAAGCCAAGGTAACGGAAAGTTTCAATCTGCTCTACCCTCTTAGCTTTACTGTTGCCTTTATAGCATTCGAATTCGAACTTAAAAGTGGAATGTTTGAATTTCAATTGCAGATCCTGTTCAAAGTTAGACTGACGCTGAATATCTTTATGCAGCTCATCGAGCGTTGTACCC tpg|BK006948.2|:84989-86381 7X32=64S 1=175S 
 tpg|BK006948.2| 821940 + tpg|BK006948.2| 821678 - INS ATTAAGATATAATGACACTATATCCTTAAACGGAAAGCATACATTCAGTGAGAAATGGGGTGTCAACAATATATCATTGTTAAAATATAATTCAGAATTGGTAGCTACGAAAGATATTCAATAGATGTAAATATTCATGACATTATCTATGC tpg|BK006948.2|:821360-822258 7X88=26S 3S1=18S 
 tpg|BK006939.2| 465763 + tpg|BK006939.2| 465885 - INS CCTCTGCATTTTTCAGCAAAGCAAGCTCCCTTTCCAGCTTGAATCTATGTTCACGCTCATCCGACAATTCTTTTTCATACTTTCTTTGTGTACTCGTAAGCACTTTTTTAAACTCACTTGTCATTATTGAAAGTGAACGTGATCCAGAACCGCTTGTGGGGCTTCCTACAGAGGAAGGTGAACTTGGATCCCAAGTCACCGGCGAACTCGCTGGTGATGAC tpg|BK006939.2|:465307-466341 7X84=26S 2S1=18S 
 tpg|BK006939.2| 66702 + tpg|BK006939.2| 67093 - INS AACAAAACAGAAAAAAGAAAAAACCCATTTGAATATAAAAATCATTGATGCAAAAGAAAGCCGTTAAATCTACAATGCCACGAAATTATTGTAATGTATGAAAAAAAGGAAGAGGGTAGCAATCCTAAAACAAAAACCCTAACAATACACATGATGCAACTGGAACGCATCAGTATTTGTAGGTTTTTATTTCGCGGATAGCGTTGCCATCAACGTCGACCTCGGTGGATTCACTAC tpg|BK006939.2|:66214-67581 7X122=55S 1=101S 
 tpg|BK006948.2| 550589 + tpg|BK006948.2| 551101 - INS GCTTAATAATAAGATAGAAAAATGCCTGCTACTTTACATGATTCTACGAAAATCCTTTCTCTAAATACTGGAGCCCAAATCCCTCAAATAGGTTTAGGTACGTGGCAGTCGAAAGAGAACGATGCTTATAAGGCTGTTTTAACCGCTTTGAAAGATGGCTACCGACACATTGATACTGCTGCTATTTACCGTAATGAAGACCAAGTCGGTCAAGCCATCAAGGATTCAGGTGTTCCTCGGGAAGAAATCTTTGTTACTACAAAGTTATGGTGTACACAACACCACGAACCTGAAG tpg|BK006948.2|:549985-551705 7X138= 277=7X 
 tpg|BK006939.2| 530414 + tpg|BK006939.2| 530175 - INS GTAACAATAAGATATCTCCTCCATTAACTTCTGCGGTTACTTCAGCTTCTGTATCGTCAATTTCAATGAAGGATGATTCAACTAAGTCATTCAAACAAGTTTCAACTAAATTACTCAAAAAAACTGAAATTCCATGTGGAGACGTATCCCTTACGCCATAATAGCTTGGATTCACATGGATACGACGATAGAAATACGAATATGTAAACCAGTCAACACAATCTTGTTTGCTTTGTATAATAGAATTTGCT tpg|BK006939.2|:529659-530930 7X171= 236=7X 
 tpg|BK006939.2| 180285 + tpg|BK006939.2| 180883 - INS ATCCCCCTCCATTTTACAATGAAATGTTAGAAAACACGGTTCCAGAAATTCAAAGGCAGAATCTTTCTCATACTATTTTGATGCTAAAGGCCATGGGAATTAATGATTTATTGAAATTTGACTTCATGGATCCCCCTCCCAAAAATTTAATGCTTAACGCACTGACAGAATTATACCACCTGCAGTCACTAGATGACGAGGGAAAACTAACAAATTTAGGTAAAGAGATGTCCTTATTTCCAATGGATCCCACTCTATCACGCTCTTTATTGTCATCTGTTGATAATCAGTGCTCGGATGAAATTGTTACTATAATCTCAATGTTGTCAGTAC tpg|BK006939.2|:179605-181563 16S157= 93=81S 
 tpg|BK006948.2| 147604 + tpg|BK006948.2| 147784 - INS AGATCAAGTAGGCAAGTATGAATTAGTTGAACATAAATTAAAGGAGTTTATGAAGTTGGATGCCTCCGCTATTAAAGCCCTTAATTTATTCCCACAAGGACCACAAAATCCATTTGGTAGCAACAATTTAGCTGTATCTGGATTTACGAGTGCTGGTAATTCTGGTAAAGTAACTTCTCTTTTCCAGTTACTGAATCATTGCAAAACAAATGCTGGTGTTCGGCTTTTAAATGAATGGTTGAAGCAACCACTGACCAATATTGACG tpg|BK006948.2|:147058-148330 7X116=17S 10S1=264S 
 tpg|BK006939.2| 69597 + tpg|BK006939.2| 69838 - INS GGGCAATAGCGCTGAGAGATTGCTGTTTCTAAGAAGCGTGGGCGAACGCAATGAAATTGGCTTTCCCTCTAGATTCAAGTCGGCGCATTACAAGAAACCGACAAGAAGACACAAATCAGCGAGGCAGTTGATCTCGGACGAAAACAAGCGGATCAACGCCTTGTTGACCAAGGCTAACAAAGCTGCAGAGAGTTCTACTGCTGCTAGGCGACTTGTGCCCAAAGCGACGTACTTTAGCGTGGAAGCGCCACCGTCTATCAGGCCTGCCAAGAAGTACTGCGATGTTACTGGGTTGAAGGGCTTCTACAAGTCGCCTACGAACAACATTCGGTATCACAACGCAGAAATC tpg|BK006939.2|:68885-70550 7X268= 328=7X 
 tpg|BK006939.2| 308820 + tpg|BK006939.2| 308680 - INS ATATATTGTACCAGGCCAATTTTTCACCTGAATCTGTAACAATTCATAAGGTTTCTCTTGATCATGATATGTTAGCAGAATTTTTCTTATGAGAATTGCGTCATCATCATCATCATCATCATCATCACAAGCAGCAGCAGTAACAGCAATATTACTATTGTTATTGTTATTATTATTGTTGTCATTATCATTATCATTATCAGTACTATAG tpg|BK006939.2|:308244-309256 7X240= 198=7X 
 tpg|BK006948.2| 394666 + tpg|BK006948.2| 394978 - INS TGTAGCCATCATTGAAAAGCAAGCGCTAAGAATGGCGCGGCGCCTATTTCTTGGTTCCAAACCATCAATAGAAATTGTGTGAGTAATGGTGGTCGCACTTGGACCTTCAGGAATCATATCACTATCTTCAACACCTTTACTTTCACTGGTATATATAGAGTTTTCGAAGGGTATCAGATTGATAAATTTTGCCTTGTGCTCCTCCTTGATTA tpg|BK006948.2|:394228-395416 282S21= 106=7X 
 tpg|BK006939.2| 374253 + tpg|BK006939.2| 374951 - INS CTTACGTAATAAAATTGAAATCATTTTCATTTGTATCCAGTAAATTGAGATCGTAATCCGGTCCTTGGTCTTCAACCATACCAATATTCCCAAACTTCAAGTTCTGAGAGTGTACATTCTGATTTTCATTAGTACTGGTTTGCTGAGGACCCAAAGTTGTACCCACATTGGATGAGGGCTGAATTAATGTGTTATCATT tpg|BK006939.2|:373841-375363 13S135=33S 18S7=7X 
 tpg|BK006939.2| 150033 + tpg|BK006939.2| 150085 - INS TCCGCCATTTTTATTTTTTATAGGTTTCTGGCAACCATGATTCATCAACTTTTTTGACAGTGGCACTCTTCTTGGAAGGTCTTTGATTTGTTTTAGACTTCATGTAGTAATAACTTACACCTCCGATGATGGCTAGAAAGATGACCTGAACTGATAAAAATTGTGGGTTGAAAAAGGAAATAGG tpg|BK006939.2|:149651-150467 7X92= 148S4=7X 
 tpg|BK006939.2| 500765 + tpg|BK006939.2| 500939 - INS TCGTACTGTACTGCCGCGTTCAAACTTAAAAGAAGTTACAGCAGGTGCAAATTCCACCCCCAAAAACCTAGCAGCTTTAATTGCCACAGGATTCTCAACCAAACAACAGTTACCAGGTATCATCGTTGGTGCAAAAACTTCGATGTTTCCAAATGTATTCTTGGTTATTTCACCGCTCGCACTGGCTAATGGAGGGATGTATAATTCTGTGTCTTCAAAGCTATATAA tpg|BK006939.2|:500295-501409 7X6=187S 114=7X 
 tpg|BK006939.2| 287348 + tpg|BK006939.2| 287933 - INS CACATTTGCGTATTGAAAATGAAAAAAAAATAATTCATTTGAAGCACTACTATTACAAAATTTATTCCAGCCCAACATTCAGTTTGGAAGCATCAAACGGCCTTCGACCATATGAAGATATTCCAGTAAATATGGTCTCCAAGCAGTTCAACTACTTTTCATGAATGTAGCATTTTCAAGGCACCTCTAACAATAAAAAAAACGACACCAGCAGGATTTGAACCAGCGCGGGCAG tpg|BK006939.2|:286864-288417 8X176=28S 1=202S 
 tpg|BK006939.2| 100911 + tpg|BK006939.2| 101133 - INS GTGTTGAGACCAAGATTATTCGTCGGTATGATTTTGATTTTGATTTTTGCTGAAGTTTTGGGTCTATACGGTTTGATTGTTGCTTTGTTGTTGAACTCCAGGGCTACTCAAGATGTTGTCTGTTAAGGCAGCTTCTGAATCACTAAAGCAGGAATAGAGTATACAAAAGAATCTTTTTGTGAGAAACTATGAAAACTATCAAAATTTTTCATCTTAGAGATTGTTTATAGCCCCTATTCTTACT tpg|BK006939.2|:100409-101635 7X8=151S 229=7X 
 tpg|BK006948.2| 634404 + tpg|BK006948.2| 635068 - INS ATATGGACAGCCAAGCATCCAGAACTACTAGAAGTTCAATTGCAATATATTTTTAACGGTTTTCAACTGCATGAGGGTTCATCGGATATGCAAAGTATAATCACTGCATCATCACATGCATTAATGTTCTTCTGTTCGGACTGCTCTAAACTATTAGTTGGGTATATTGA tpg|BK006948.2|:634050-635422 7X1=1I88=37S 1=363S 
 tpg|BK006939.2| 546013 + tpg|BK006939.2| 546160 - INS GATGAAGGGTGTAATAATTTGTAGTTCATTATTGCAATTATATATCTATATCTATATATGTATATAACATTAACATGTGCATGTACACACGTAATCGCGCGTGTACATGTCTATATGTGTTACTTGAACTATACTGTTTTGACGTGTATGTTTATTTATCTCTCTTCTGATTCCTCCACCCCTTCCTTACTCAACCGGGTAAATGTCGCATCATGACTCCCGACAATAATCC tpg|BK006939.2|:545535-546638 13S169=28S 24S5=7X 
 tpg|BK006948.2| 570872 + tpg|BK006948.2| 571504 - INS ATTGTAGGCAACACCTTTGTATGTTTCGTTTTAGCTGATGCAACTTGTAAGTTCGCAACCTGCAACTTACACTTCACCAGCTCCACGGGTGTCAAAACTAAACTAGCACATGAACCCGCTACTCCACCAGAGATCAGGATTTGCCCCAACGGGGAAACGTTTGTATGTTTTTCTACA tpg|BK006948.2|:570504-571872 7X6=82S 76S11=1X1=7X 
 tpg|BK006939.2| 152433 + tpg|BK006939.2| 152138 - INS TTGTTGAGCTTAAGACAGTAGTATAAAGTCTTGTTTAGTGCAAGCCACTGTTGGCGTTTCAACTAAACTATTCCTTAAAAATAAAGTACAATGTTACTGCTAAACAATGTTGAAGGTGAGCTTAAGACAGTAAATCAAGGAAATGCGGTATAATTCCTGCTGACAAAGCCGCACATAAATAGCAGTTGTTAGCTATAAGGAGATTTTTAGCTACGAACATGG tpg|BK006939.2|:151680-152891 7X3=329S 195=7X 
 tpg|BK006948.2| 440163 + tpg|BK006948.2| 440581 - INS ATATATATGGTGATACCCAAAATTAGCTTGGACAAAGTTTCATTGAATTGAAGCCGTTTGTCATTAATATGCACGTTGCGATACACTTCCGTTTTCGTTCCGATCTTCCTTTGTTGAGATTGTTGTATTATTATATCAATACTACCTTCCTTTGATACGGAGGCCCTTGTC tpg|BK006948.2|:439807-440937 19S157= 150=7X 
 tpg|BK006939.2| 155502 + tpg|BK006939.2| 155378 - INS CATGGTGCTAAAGCCATATAGTTATAACCACAGAACCACTCACGGCGAATTAATAACTCTAGATGAGGAGCAGCGCCTACATATTGATGCTGTCAACACTGTTTGGTCACATGCTAATAAAGATAACACCAGATCATTCACTGAAGAAGAGATCAAGGAATTAGAAAATTCTAGACACGAACAAAGCTAGAATGCATTAACCAGTGTTTTTTCTAACTGTTTATGGTACTAGCCTTTGTGAACATGTATAGT tpg|BK006939.2|:154860-156020 7X259=1X28= 126=7X 
 tpg|BK006939.2| 163941 + tpg|BK006939.2| 164056 - INS GTCTAGTTTTCCTACAATCCCATTAAGAGCTTCTTCTGGTGCAGTCAACGGAACTTCTTTCAACAGAAAGCTAAGCCAAACCACTACTGCAAGTGCACTGCTAGAGTCGCTGAAAACTTACTCTAATAACAGCAAT tpg|BK006939.2|:163655-164342 7X4=64S 64S4=7X 
 tpg|BK006939.2| 324893 + tpg|BK006939.2| 324311 - INS GAGAACACTGGTCTTCTGAAATTAGGCCTTGTTTGATTTGGTGGTTTCTTTTACGAATATTTTTCTCCTTATCCAGTTGTTTCTGTACTCTTAATTTTCTTTCATCAATAACGTTTTGAGTCTTTTTACGCAAAAAGGAACGCAAACCCGAATTCTTACCTTTCACATCAGGTTTTACATCTGGAATGTCGCTGTTGGTTTTGGCTTTATTATTAGCATCCATTGTAGTTTGCGCCAAATCCTTAGCG tpg|BK006939.2|:323801-325403 7X4=163S 233=7X 
 tpg|BK006948.2| 414360 + tpg|BK006948.2| 414839 - INS CTGCTTCATGACCTTCACTTTTCAATTTCCCATATAAAACGTTTGCGGTTTTTTTGGTTGCAACAAAAATAATGGAAGATCCAATTGTCATTAAACCATATAGCTCAGTTAAAACATCAAACTTATCTGCTTCGTTTTTGCAGTCCATGTATAGTTGTTTGATGGCATCAACATTAACTTCATTTGTTTGTAATTCTAAAGTATTAGCATTTGGAACGATCTTCTTTGCGTACTGCCTAACTGCATCGGCAAAAGTAGCACTAAACAAAACAAGTTGAGTATCCTTGGGTAAAAATCTCTTAACACGAATACACTGGTCACCTAGACCCTGCTGATCCAACATGTTATCGGCTTCATCCAAAACAAAAATTTTAATTTTCTGTAGCTGCATCAATTTTCTACGCATTAGGTCAAGAACAGTGCC tpg|BK006948.2|:413498-415701 13S17= 212=7X 
 tpg|BK006939.2| 206144 + tpg|BK006939.2| 206202 - INS TGTTGGTACTAAAGTTGATCCTACCTTGTGTAGAGCTGATCGTCTTGTCGGTCAAGTCGTCGGTGCTAAGGGTCATTTGCCAAACATTTATACTGATATCGAAATCAACTACTTTTTGCTACGTCGTCTATTAGGTGTCAAAACAGATGGTCAAAAG tpg|BK006939.2|:205816-206530 7X90=27S 7S1=156S 
 tpg|BK006948.2| 509067 + tpg|BK006948.2| 509518 - INS TTCCTCCTTCTTGTTTACCAAAAGAAAATATTGGAGCAGTTGATTTTGGAGGCGCGTCTGATTCTGTATGATTTTCACTTTTTTCGGATGTCTTTCCAAATTTAAAAGGTTGACTGGCAGAAGTAACGGTATCTGATTTACCACCAAAATTGAATAAAGTTGTGGAAGGGACAGTATTGTCGAC tpg|BK006948.2|:508685-509900 13S85=47S 39S7=7X 
 tpg|BK006948.2| 335477 + tpg|BK006948.2| 335037 - INS GTTACAAAGTGTGTAACAATATATCGTACCGTATTCCAGTGTCCTCCGTGACATAGTCAGAGAGAACATAAAAAAGTAATCCGGCAAAGATGTTTGAAATTGGCAGTTGTTTCCTGTTTTGGTGAAAGCTGTCTGAAATAAGTACTCTCTTTCTCTTTTTCCGTATCAATCCAAGCTGTGACCTTTCCGCTTGATAGCTGGGGTTAGATTTAACCGTCCTACTTTCGTATAAGTCGTTAAGTGTGTAACAA tpg|BK006948.2|:334521-335993 7X193= 13S223=7X 
 tpg|BK006939.2| 348177 + tpg|BK006939.2| 348642 - INS TTTATGGCCTCATGAGTTGGATGTGGAAAATTCTTGACGTTCCGCTGATATTTTGTGTTGGGGTTGTTTTTGGGACCATGAGATTGCCATGAACCGATCAATCTTGTCTCATCTTCAAGTATCTCTTCACCACTTCATCCTTCTTGATGATGTATACTACAGCTCCCCAGCCTGATAGAGCGTCACGGTCAGCAGCATTCAGTAGGGCCTGACTTATAGTTTCGAAAAGATCTTCTGGCTCTAGATTAGGTTCGTACAGGGACTCACACATACCGAACAGTTGGTCGGATGCAGTACCGC tpg|BK006939.2|:347563-349256 7X24=1X162= 282=7X 
 tpg|BK006948.2| 862654 + tpg|BK006948.2| 862642 - INS GATCCTGATCCTGACCCTATTCAATGAAGTGTTGCATCCGTTTTATGTCTTTCAAGTATTTTCGATAATTTTGTGGGGCATTGATGAATACTACTACTACGC tpg|BK006948.2|:862424-862872 7X6=79S 5S85=7X 
 tpg|BK006939.2| 412072 + tpg|BK006939.2| 412347 - INS GGTTACCATGAAATGATTAATCATTGTTGTTTTTACAGCAACATGGAAAGCAGCAAAGAAAATGCAGGAAAACGTGAAGTGCTTTTTTTGATGATTACGCAAAGTTCTTTTCAAGTTCGCCATAAGAGGAGGTTTTCCTTTTCAAAAGGAGCATGATACCAATAATTTATATTGCCTTACGC tpg|BK006939.2|:411694-412725 7X8=83S 87S4=7X 
 tpg|BK006948.2| 583969 + tpg|BK006948.2| 584180 - INS TCGTGCCATGCTTGATGGCTTCTTGAACGACAGAAGGCGACGAACATTTTTTCACCTTGAATTCTGTTCCCAACGTATTACTTTGTATCCATGACCATGCACCGTTTCTGCTTCTGATAAAGTATGAATATGGCGATAGTGCTGCCATTGTGAGGATGTAGGGATTTTCGATCAGTCCCAATTGCTTTGCAGTGTTGATTATGTGTGTCTCTGGATGTGAAAGGTTCCATTCTCCATGCAGTTTGGACGCCAAGTCCTTATATTCCTCCATTTTAGCGGCTCTCGCAGAATTTAATGT tpg|BK006948.2|:583359-584790 7X234=26S 1=52S 
 tpg|BK006948.2| 619753 + tpg|BK006948.2| 619896 - INS GAACTCAATGGAAAACAACACCACACGTATGATCTTACTAATAAAAGCACATGAACGTTCCTCAGCGCGAACGTTCGCATTCTGCGCCTTCGAGCACAGGATAAGTTGCAGGAAGCCATCACATCTATGCAACGATTATCACGACACAACCTTGCCGCCGAGCA tpg|BK006948.2|:619411-620238 7X6=76S 77S5=7X 
 tpg|BK006939.2| 442941 + tpg|BK006939.2| 442275 - INS GTGCCCTGTGCGGCAAGGTAGTTCTGGGTCCTTAGGGGCTCCACCTTCACCGCTGTTAGGGGAGTTTTATCCAGCGTCAGCAAAGGTGACCCGTGATGGAGGCGGCCGGGATAGCACATATCAGTCGGATAATTGTGCAAGTTGATCGCTTCGGCGGTTTAATTTGGCGGTGCCATCAGGATTTACTCGCACATTGTGGCCGTTCCCTCGGGGATGGAG tpg|BK006939.2|:441823-443393 7X4=154S 110=7X 
 tpg|BK006948.2| 175469 + tpg|BK006948.2| 175733 - INS GCTACTATTCCTAACGCTATCTTACTTGATTCTATGAGGATGATCTATAAGAAGTGGCATACTTACACACACAGTAAAAGTTTAGAAAAACAAGAACGGAACGACTTCAGAAATTTCGCGGGTATTTTAGCCTCTTTGTCGGGTATCCTATTCATCAATAAAAAG tpg|BK006948.2|:175125-176077 7X4=78S 76S7=7X 
 tpg|BK006939.2| 449685 + tpg|BK006939.2| 450078 - INS GAACCAAAACTCTGAAGCAACACTTTCGTATATGGATGGCCCTTCAGAGAAACCAATAGGTATGTAAAGAATTGCTACGTGGTGACTCAAAGTGAATTATAGCAAAGTTATAAAAGCGCTACATTGTAGAAAATTGAGAACCACATTTTGACA tpg|BK006939.2|:449365-450398 7X115=18S 1=198S 
 tpg|BK006948.2| 549171 + tpg|BK006948.2| 549750 - INS TTATAATCTCATTTTCCACAGTCGCCCTATTTGCTTTATCCTTTGATGTTTTCGCTCTGCTGAATGATAATTCATCAGTTTTTATTTTGTGACTATACTTCTCTAAGAGCTGATTATTAATATGGTCCGAGGCACCTTGCGACACAGACAATGAATCAAATTTATCTTCCAAGGACATGACCTTCGAAAAATAACGGAGTTTGAATCTCTAAATCTGTTTTAACTTCTTTTTACTATTATTTTTAGTCTTAGTATCTCATCTCATCTCAATTTCTATATTCCACTATAAAATTTTTCACTCTTTCTGCG tpg|BK006948.2|:548539-550382 7X8=11S 166=1X123=5X2S 
 tpg|BK006939.2| 457738 + tpg|BK006939.2| 458191 - INS GACAAACACAATAGCTTCATGGAAGGCTGCTTTTTTAAGCATTTAGGACATGACCATTGTTCATCGACACCTAACCTTTCGCATTTGGTGAATTCCCGGAAACAGTCTAATATGTTACAAGTTTTAACGCGTGGGACAGGAACAGAAAGAACAGAGAATGTTTGGTAAGTTGTGGAGGTATGTTCACAAACTTGACATTGTAGCCTAGATGCGTACTGTCCTTGGAAAAGGTCAATTATCGCACTGAAGTCGGTAAGCAAAAATCTTTCCCACTCGAGAGCACTAGCTTTGCGTATGGACATTTTTTCTCTCATTCGTTCTTCCTCATCTGATAACTGTTTAAGATGCTTTTTGCTGCCGTTTTGGTTCAAATC tpg|BK006939.2|:456976-458953 8X13= 351=7X 
 tpg|BK006939.2| 39020 + tpg|BK006939.2| 38736 - INS TTGAGATCTACTTGATGGTATTCGGCAGTGATTTTGTCCCTAACCTTTTTCTTAATAGAGCAGCTTTAGGTGTTAGATCATTTAATGACCTCGGAGAACTGTTCCTAGAATTACTCCTGGAACTACTAGCACTGTTGCTAGTGGTATTATTTGCTGTGCTTGAATCAAAAATCCTCAATTTTTTCATAAATTGGCCGTCAAAGCCAGTATTACGAGAGCCGTTGCTATTGC tpg|BK006939.2|:38260-39496 7X6=4S 25=1X173=1X17=7X 
 tpg|BK006939.2| 239476 + tpg|BK006939.2| 239840 - INS GGAAAACATTATTCGAGGAG tpg|BK006939.2|:239422-239894 7X5=5S 10=7X 
 tpg|BK006948.2| 229269 + tpg|BK006948.2| 229649 - INS AGGAATTTGGTATGAGGATCAGAAGGAGGTTACACGGATACAATCGAGTTCTGATTCCGAAGATCGTTCACTTTCGTATTCCGGCTCCAGCGATGTCAAGGATAACAATGACGATAACACGGAAGAATTAGATGACCCACAACCGAAAAGGCAGAAACGCTTCCGTGTAGTTCTAGG tpg|BK006948.2|:228901-230017 7X197=1X12= 155=7X 
 tpg|BK006948.2| 610743 + tpg|BK006948.2| 610815 - INS ATATCTAAAATAGTGAACAAAGGCCCGTAAACCAATAATAGGGGGCCGTAACTCCTAGCAGCAAATTTTGATTTAAATTCCCATGGGATGGTACCTTTGACCTTCATGAACTGCATAGCCAAAATCTCGATGCATTGGAAATGTTCATCTGGATGAATATACGACGGGCCTAGGC tpg|BK006948.2|:610379-611179 7X2=1I18=66S 3S1=175S 
 tpg|BK006948.2| 311169 + tpg|BK006948.2| 311382 - INS GGGGCGGAGGACGGTACTTCTTTACTTTACCCTGACTAACATTTGATTTTGGAGTAGAGCGGTCTTCAGAGTCGGGACTTAAATTGTATGATGTATAATTGAATGGATTAGTGCTGTCTGTAAACTTTCCCAGTATTTGGGTAGCACCAGGTTCCCTTGGAGTACTGGACAAGGAATCATATAT tpg|BK006948.2|:310787-311764 7X6=199S 92=7X 
 tpg|BK006939.2| 342944 + tpg|BK006939.2| 343570 - INS CATTCACAGTTCTCAATTGAGCAGAACGAGCTATGACTACCACAGTTTTGCGACCGGGAGATAGAGCGAAAGAGCTGCCATGACTGCGATGACTCTAGCGAAAAATATTGGCCTTTTGCACGTTCGCGACTAAACGAGTTCGATAGTAGTCCCGTTTCTGGTTTTTTCCCTTTACCGGCCCACATTTTTTCACCTGACTCCGGTCCTGACGTACGACTCTGTTTGTAAGTCACGTGAAATATTTCCTGTG tpg|BK006939.2|:342430-344084 7X5=224S 125=7X 
 tpg|BK006948.2| 346034 + tpg|BK006948.2| 345358 - INS CTCCTCTCCTTACAACTCCACAACCACCACCACCCCAGCTAGTTCTGCTTCCAGCGTTATTATCTCAACCAGAAACGGTACCACTGTTACTGAAACTGACAACACTCTTGTCACCAAAGAAACCACTGTCTGTGACTACTCTTCAACATCTGCCGTTCCAGCTTCCACCACCGGTTACAACAATTCTACTAAGGTT tpg|BK006948.2|:344952-346440 7X5=168S 98=7X 
 tpg|BK006948.2| 640779 + tpg|BK006948.2| 641153 - INS CATTCGCCCATAATTGTTTATATTTTTCAATGAACCCCCAATTACTA tpg|BK006948.2|:640671-641261 7X5=18S 20S4=7X 
 tpg|BK006939.2| 317561 + tpg|BK006939.2| 317976 - INS GTTCAATAGTAATAACTTGTCCAACCTTTAATGGTTCGTACCTGGAAACTTTAGGCACATCGTGAACATCTAGACCTAAATTGTGTCCAATATAGTGCGGATACAATTTTTCAACATTCCAACCGGAGACTTTATCTATGCCCAAGTTTTTCAATTCCTGTTTCATGAGTGTGAT tpg|BK006939.2|:317197-318340 7X5=82S 84S4=7X 
 tpg|BK006939.2| 565760 + tpg|BK006939.2| 565966 - INS CGCCAACACTATAACACTCACTGATCATGTGCTCAATGGGCAAACATTGTCTAATGG tpg|BK006939.2|:565632-566094 7X7=55S 29=7X 
 tpg|BK006939.2| 271087 + tpg|BK006939.2| 270459 - INS CCATAATTCTAAAAGACGCTATTAAGACTTGCCCTTAATCTCTTTCGGCAGCAATGGCTGCCATTTCCATGTCAACGCCTAATGGCAATGCTGCAACAGCAACGCATGATCTGGCAGGTTTGTGAGTATTGAAGTACTTGGCGTAAACGGAGTTAAACTCAGCAAAGTGATTGATATCTGCCAAGAAAATGTTAACTTTTACGACCCTGTCC tpg|BK006939.2|:270021-271525 7X4=265S 106=7X 
 tpg|BK006939.2| 141579 + tpg|BK006939.2| 141269 - INS CAGGTTATGTG tpg|BK006939.2|:141233-141615 7X3=2S 6=7X 
 tpg|BK006939.2| 154223 + tpg|BK006939.2| 154573 - INS GTGTTACTGTGTATTAAATGTTGGCACTCCGGAGATTTATATTAAACCAAAGGTCTTTGAGATCGTGTACCATACCGATTCTAGTCGGAGCCTTGATCATTATTCTCGTGCTATTCCAACTAGTTACCCACCGAAATGATGCGCTTATACGATCAAGCAAT tpg|BK006939.2|:153887-154909 7X4=76S 77S4=7X 
 tpg|BK006948.2| 145227 + tpg|BK006948.2| 145683 - INS CCTTCCATCGATTATGAACCAATACAATGTCGATACGCAAGCAACCGCTATAATGAGCGATATGCAAAAGCAATACGACTCGCAACAGATGACATCACCATTTGTAAACGAAGACTTGCATTTCGATCCAAATGGTGAAGTTTCACACGTAATAAAAGCAATTTTTAAAGA tpg|BK006948.2|:144871-146039 12S12=1X107=24S 15S7=7X 
 tpg|BK006939.2| 220030 + tpg|BK006939.2| 219798 - INS GATGATGTCCTTACGTTTGAC tpg|BK006939.2|:219742-220086 7X10= 6S5=7X 
 tpg|BK006948.2| 959539 + tpg|BK006948.2| 959849 - INS CCGTCCTAATCACTTGTGGGTTTGTAACCTGTTTTTTGTGTTTCTTGATGAACCTTGCGGTTTCGCGGTTCTCATTGGCTCTTTTTACTTGTGACATAATCCACGTTTGTCTCTTATCTTTCTGATATTATTATATATAAGCAAAAAAACGAGGGAGTGTATAACGAT tpg|BK006948.2|:959189-960199 23S68= 30=61S 
 tpg|BK006939.2| 2080 + tpg|BK006939.2| 1607 - INS TCCGTATTGTTGGAGTTGGTGCTAGCAGTGGTAGTAGCACTAGTTTTGGAGTTGGTACTTTCAGTGGTAGTAGCATTAGTGTTGGAGTTGGTACTTTCAGTGATAGTAGCATTAGTGCTGGAGTTGATACTTTTAGTGGTAGTAGCACTAGTCCTGACGTTGATGCTGGCAGTGGTAGTCGCATTAGTGCTGGAGTTGGTACTTTCAGTGGTAGTAGCACTAG tpg|BK006939.2|:1147-2540 14S104= 112=7X 
 tpg|BK006948.2| 125891 + tpg|BK006948.2| 126585 - INS AAATATATAAGTAATAATGTGTCAGTAAAAAAGAACAAATACATCACGAAGACAGAAATACGGACAAGAACCGCAGAAGACATTAAAGTCAAAACATGAAGCTTAATTCAACTCGTGTAAGT tpg|BK006948.2|:125633-126843 25S43= 18=50S 
 tpg|BK006948.2| 369918 + tpg|BK006948.2| 370327 - INS GTACACATAGTGTACACATAGTGTCCCTAAAATTCCTATTGATGAATAGATCAATTTTATTAGCAGACAATTGGGGGCAGCAACTGAATAGCAGAAGAAATTTGAGTTCAATTATTTTTTTTTCCTGTCATACATAATGGCCTATTTACAGGTACATACATATAGAG tpg|BK006948.2|:369570-370675 7X12=147S 147=7X 
 tpg|BK006939.2| 103976 + tpg|BK006939.2| 104077 - INS ATATGAACAAAAAGGTATTTCTCGGCACCATCTGAGAAACAGCTCACAATACTCTCTTTAGAATTGAGCCCATGGATAAAAAATTCTTCTTTTTTACGTAGAAAACCAGATTTTGCCTCAAGTATCGAAATCCTGAGCTTGGAGTTCTGTACGGGA tpg|BK006939.2|:103650-104403 7X1=1X3=1I19=53S 71S7=7X 
 tpg|BK006939.2| 61538 + tpg|BK006939.2| 61410 - INS TTCATCATGGAACTATACT tpg|BK006939.2|:61358-61590 7X3=6S 7S3=7X 
 tpg|BK006948.2| 283944 + tpg|BK006948.2| 284156 - INS TTTGTATCCTGAAATCTGAAAATGTGTCCCTTTCAAGATCTTTATCAAAAGAATCCATTTGAGGAATAGAGTCTCTGATGTCGTCTGCATTTGGTAGTAACTCGATATACTGTACCAAGCTCTTGGTTATTATATTGGACTCCACTTCCTTAGTGGCAGCTTCTCTATTCAAACGATCGTTGGTAACAAGAACGACGTTTATGTCATAAGG tpg|BK006948.2|:283508-284592 7X7=98S 100S6=7X 
 tpg|BK006948.2| 1060767 + tpg|BK006948.2| 1061183 - INS CTGCTGTTGGTGTATTTGGCACCAGGTTCTTTAGCAAAACCAGCATCAACTAAGAAAAGAACGCAATGGGACCAGATAGCAATTGATGCTTGTGCTAAAGAATTGGAATCACACAAATTTGACACGGATGTGAAGGGTCGGCACGCTACTCTTTGCACTTATGAACCAGCACTAGGGTCTTGGTTACATTGCGCGAAGGATGTTCTCGACAGTAGGAAGAAAAGTAAAAAAATATTCGAAAAAACGTTTAGCAAAATTAATCAGTATTGCCACGATTATCACAAAGATGAGGTCGTCAGCAATGAGGAGTATTATCGAATTTTTGCCAATGCATCCC tpg|BK006948.2|:1060079-1061871 7X287=28S 5S1=62S 
 tpg|BK006948.2| 789464 + tpg|BK006948.2| 789370 - INS ACTGGAAATATCGTAAAAGAATATAGATACGCATAATTTTCTTGATACAATAGGCGTAATTTCTAGAACCTCTCCAAAATTCTGAAAATCTTTTTCTAATTCTTGAATATCAATGTTTTCTAAAGTTTGCCCTTTATTCAGATTTGATTTGTTAGGCATT tpg|BK006948.2|:789036-789798 7X5=75S 76S4=7X 
 tpg|BK006948.2| 720842 + tpg|BK006948.2| 720815 - INS AATTGGTCAACAAGTTTAATCTGTGCTTGTCCACCAGCTCTGTCGTAACCTTCAGTTCATCGACTATCTGAAGAAATTTACTAGGAATAGTGCCATGGTACAGCAACCGAGAATGGCAATTTCTACTCGGGTTCAGCAACGCTGCATAAACG tpg|BK006948.2|:720497-721160 7X4=72S 69S7=7X 
 tpg|BK006948.2| 806448 + tpg|BK006948.2| 806823 - INS ATACTCGCTGGAACTTGAGCCCCCTCTCCGAAATACACATTGAGGACATGATAAATGAACCGTCTGGACTATGTCCAGGAAGTTCCAAAAAGAAACCACTACTGATTGCAAGGTTTCCCAAGGGTTGCCAAGAATCACCAAGGGTATATGTACTGCAA tpg|BK006948.2|:806118-807153 7X7=72S 74S5=7X 
 tpg|BK006948.2| 1048475 + tpg|BK006948.2| 1048520 - INS AAATTGATGAACACCTAATGTAGTCATTTCCTTTCTCTCTTTGCTAGTAGATTTTAAAAAGGTTTCTTGCTGTATTTTTTTATACTTTTATAGACGCCGCTTTCCAAAGTTCATCTAAAATAAGTCGCTACAATGATTTGATCTTGATTCGGTGCTTCAGGAGCCTGCTTGCTTCTTTGCAGCTTCGGCAATTTGGAACCTTGTGTGCATATCCTCGTTTGTAAGCCCAGAAG tpg|BK006948.2|:1047995-1049000 7X52=1X97=1X27= 219=7X 
 tpg|BK006948.2| 673463 + tpg|BK006948.2| 673600 - INS CTCCTTATATTTATTACTACGCAGATTTCGAGTAGTTGTCACATCAAACAGAATAAAAGGGGTATTGTAAATTTACTGACTTTTCCATCAATCCCGTATGAATGGATGGCTTACATATCTTGGAACGCAGACTTCGAAATTAAGTATTTAGGAGTGAGAATGTGCGTTAGCATTTTGTCTCATATCTAAATATTCAAGTTTAACTTGTATTATTTGTCCTCAGTACAAGAGGTGTACGGCTTTTGAAAGTCCACTCCCCCATTTTTATCC tpg|BK006948.2|:672909-674154 7X13=9S 135=7X 
 tpg|BK006948.2| 1018755 + tpg|BK006948.2| 1018906 - INS TACGACACAGGCAACGGTGATTTAGCTATCGGAACCCATTATAAATTGTGAGGAAGCTTACCAACTCATAAGTGGAATAAAGACACAGGCAACACTTTTCAGAAGCAATGTCAGCAATGATTCAGAAAAGTGACCCCATCAGGGTCGAAATCTGAGTGCTCAGATTATCTCTTCAAAGGGTAAATTACGGGTAGGACTACATATACAGAGAACTTCTGGGACCTGGGAAATACTGTTCTTTCTAGTGTGTATACATGGGAATAGCTGCATATTTCCAGAC tpg|BK006948.2|:1018181-1019480 13S153= 263=7X 
 tpg|BK006948.2| 363226 + tpg|BK006948.2| 362821 - INS TTTCTGTATTTTCGTTGCTAATAGGGAATTTAAGATGTCTATGAATCTGTTCAGTAATATTTTGAAACACGTTGAGCAGTTACTTAACTCAAGTAATACGAAATGGGAAAAATGCAAAATAATGCTTAAAACCGAAGTTGAAGAAAAACGATCCAAAAGTGGCCGCTTCTTTAACGAACCGGTGCTAAATATTGTAGCCCTGCCGTTGTCACCTGAG tpg|BK006948.2|:362373-363674 7X265=14S 3S201=7X 
 tpg|BK006948.2| 715844 + tpg|BK006948.2| 716477 - INS TCGTCCAGATGCGTCTTTTTCCCGAAGTCCCTGTTAACTGACTGGTTGCATTTTCAACCTCAGTTGAATTTCCAACTGGTACCCTAACGCTAGCGTTATCTGAATCAGTATTCAATGCATTGGATCTTATTGGCCGAGTTGCGCTCGTTCCACACCTAATAGTGGACGAAATCCATCTTGTATTTCTCCCAACAAATAGTACTCCAACAGATCGTCTATACATTATTGTGGCTTAACAGTTCTCCTTAAAATCCACATAACTGACAAAACTGGATACTTAATGCCCATCGAGTCATATAC tpg|BK006948.2|:715230-717091 7X17= 282=7X 
 tpg|BK006948.2| 346799 + tpg|BK006948.2| 347371 - INS ATTGTGTGCTTTTTTGTCCACTCCTTTTTCCGTAAATATTACATAATTAAATAGTCACAGCTCTTACGCACCTGTTTGGCCGCACATGAGAGTTAAACGCAAACTCCGCCGAGGCGTCGTTTTTCTAGCTGCTGCTTCACGTTTTATGGAGTCATATTCTGGTCTAAAAAAATTATACTATGCAGGTAATGGATTGTTTTAAGTTTCTTGTTAACTCACATAG tpg|BK006948.2|:346339-347831 15S79=24S 108S4=7X 
 tpg|BK006948.2| 1035428 + tpg|BK006948.2| 1035984 - INS GGGTAGAGCTTGCTGTTGTTGTTGTTGTTGTTGTTGTTGTTGTTGTTGCTGTTGTATCTGCTGATGATGCGGTAATATACTGTTCTCTACCAACGACGATTCGTTGCTCGAACTGTTGTGAGCGTCTGTATTGGCAAAATGATCTTGAGTCTGTTGATAC tpg|BK006948.2|:1035094-1036318 7X12=28S 80=7X 
 tpg|BK006948.2| 710471 + tpg|BK006948.2| 710878 - INS ATGTTAAGAAAAATAATATTACATTGGATTTTTATAAGATAATACTAAACTTATTGTCTAATCTAATTAATATTAAAGGTAAAAGGGACAAATATAACTCAGAGCTAGCTTACGAAATAATTTCAGTAGGTTCCGGTGTTACTGAACTCCTTAAGCTATGGAACCGAGCCAAAGTCACTTCGGCTAATG tpg|BK006948.2|:710079-711270 7X14=80S 89S6=7X 
 tpg|BK006948.2| 835134 + tpg|BK006948.2| 835104 - INS GGTTTTTAAAAATTCTTTCTGAGCTTCCCTGCTGAACTTCTTCAAGGCTATATTTCTCTTCTTGGCACGCTTTCTTAAAATAATACCTTTATGGGTCTCTGGCATGAGCGCAATAAATGGCAAGATTAGACCGCCCGCAATCAATTGGATCCATTCAGACCAACGCCAGCCTTTGGCTTCAGT tpg|BK006948.2|:834724-835514 7X5=86S 19S14=66S 
 tpg|BK006948.2| 225707 + tpg|BK006948.2| 225530 - INS CTCTGGGATGTTGGAAAATATCCTGTAATCCGTTAACCTTTCTTTCCTCACCTAACAATTTGTAACACTCTGGGATGTTAGGAGTCAAAATATCAGCAAAAGGTGCAACCTTCTCCGTAATCAAACTAACTATATCCTTTCCAGCTAAAGAAGAACCAGAAGTAGCGACAAGAACTGGATCAACAACCAACTTAGGTCTATTTTCGCCGAGTTGCAGCAGTTTTTCGTGCAAGACTTCGATAGCAGCTGCGGTAAGCATACCGGTTTTGATAACATTACATTTCATATCCTTTAAATTGGATTCCAAAGTTTGGAAAACCACTTCTTTTGGTGTGTTATTTATGCTGTAGACTTTAACTGGAGTTTGAGCATTTAAAGCAGTGATACATGTCATGGCATAACATCTGTGTGCTGTGATAGTTTTGACATCAGCTTCGATACCGGCTCCACCACTTGGATCTGTTCCAGCAATGGATAAAACTGTTGGCAACTTTTCGTTGCAGGCTAAAGTAAGATATGGTGGAGGCGTGTTGATGCTAACTGTAGAAT tpg|BK006948.2|:224418-226819 7X6=18S 532=7X 
 tpg|BK006948.2| 219625 + tpg|BK006948.2| 219283 - INS AATATACACTAGACCAAGGCTACGAAGTTGTAGCTTTCATGGCTAATGTAGGGCAAGAAGAAGATTTCGATGCCGCCAAGGAAAAGGCCTTGAAGATCGGTGCCTGCAAGTTCGTTTGTGTGGATTGTCGTGAAGATTTTGTCAAGGATATTCTATTCCCAGCTGTACAGGTCAACGCTGTGTACGAAGACGTTTATCTGTTGGGTACCTCTTTGGCAAGACCTGTTATTGCCAAAGCCCAAATTGACGTCGCTAAACAGGAGGGCTGTTTCGCGGTCTCTCATGGTTGTACCGGTAAAGGTAATGATCAAATCAGATTCGAATTGTCATTTTACGCTCTGAAGCCAGACGTTAAGTGTATTACACCATGGAGAATGCC tpg|BK006948.2|:218511-220397 7X5=86S 190=7X 
 tpg|BK006948.2| 845238 + tpg|BK006948.2| 845812 - INS CCTCCAGTCTCGCGTAAACATTCAGAGAAGTACATGACAAAGTTTGCTGTTCTTTATATCTGTATATATTAAATAATGGGGATAGTGACACCACTTAGCCTGTAAATAAGGAATATTCGCACTATTTAGTCAAAAAATCCATCATCATCATCATTAATGTTGCC tpg|BK006948.2|:844896-846154 7X10=72S 76S6=7X 
 tpg|BK006948.2| 516368 + tpg|BK006948.2| 516359 - INS ATTACACCCTTCCTCAATTTATAAAATGTAAACAAACGAAATGTAAAATCAAACTAGCAACAATAAACTCGGCAAAAGCTCTGTTTTTAGAAATGCCTGGAAAACTATTACACAATTGTAACCGCAAACTCATCAATAGGACGAATTGTCCCACACAAATAATGAATCCCGCTAAAAACGCATTGAATGGAAAATTATCACGGATCAAGATAATGAATGTACACTGGATCACCCCTAATAATACCAAAAAGAAGCAGAATGTATCAATTAGTTTCAGTTTAGGATATTTTTCAATTTGGGCAAAATATGCCCTCTTAGAAGTCTTGAAAGTTTCTTGAAAATCTGTTAAGAC tpg|BK006948.2|:515641-517086 7X204= 176=7X 
 tpg|BK006948.2| 226456 + tpg|BK006948.2| 227096 - INS GAGTTTGAGCATTTAAAGCAGTGATACATGTCATGGCATAACATCTGTGTGCTGTGATAGTTTTGACATCAGCTTCGATACCGGCTCCACCACTTGGATCTGTTCCAGCAATGGATAAAACTGTTGGCAACTTTTCGTTGCAGGCTAAAGTAAGATATGGTGGAGGCGTGT tpg|BK006948.2|:226100-227452 7X6=79S 82S4=7X 
 tpg|BK006948.2| 249761 + tpg|BK006948.2| 250196 - INS CGTCAGGTATACTTAGGATAACTGCTTCAC tpg|BK006948.2|:249687-250270 7X5=10S 10S5=7X 
 tpg|BK006948.2| 1070860 + tpg|BK006948.2| 1070328 - INS TGTATAGGTGGAGATATATCAATTATACCTGTTATATGCTGAAAACCTTAATGATTATATTAACCTTTTTCTAGCAACTGAAAATACAGATCTGGAATATGTTTCTATATTTCCAACCTCAGCGGTTATTCGAAAAAAAAATAATTGACCCGCAGGGTGTATAGGTAGTTGATGAAAGTATCATTGTTTTTAATTTATTGTTAAAAGTCCGAAAAGCGAGAATGCATGAAAGTATTACCTTCCATTCCAGGAATAGAAGCAACACTAATTCAAAAGCCCGTTTAGGAAAGATCCGAATATTTTGACAGTAGTACGTAATGAATAACCACTCAGGTGATACTAAGACAAATTTTACAACATTTTAATGTGTTCCTGATTTGATTATGCAACACTTTTTTTGACCC tpg|BK006948.2|:1069506-1071682 7X9= 1S391=7X 
 tpg|BK006948.2| 294395 + tpg|BK006948.2| 293925 - INS AGAGAGTAACTACAACGAATGCAGTTCAGTAAACACTAGTTACAGTTTCAATGACATGTCAACTTATCTTAATTACTTCGTAAAATTCAAAGAGGAGGGTACAAAAATACTGCCTGCAAAAACCGCACAAAATGAAAACAAGTGTCAACTTAAACTTATATATAGGAACACTCCTGCATGTATCCGTAATTTACAGTTCAATGA tpg|BK006948.2|:293503-294817 7X4=231S 192=7X 
 tpg|BK006948.2| 22160 + tpg|BK006948.2| 22290 - INS CTATAATAGTATACATTTGTATCACATTTGGGTGCAATAATTTAAACAGATTTTTGCAGTTGACTCAGGACTAAGGGCAATTCTTGCCCAAACTACGGAACCCTGTTTCTGATCCGAAGGGCTTATAATCCATAGAAACCCTTACATTTGCTCACTGAAAACCCTGTGTCCTTATTTGGTATATATGATGCGAGGATTA tpg|BK006948.2|:21748-22702 7X5=94S 96S4=7X 
 tpg|BK006948.2| 344495 + tpg|BK006948.2| 343833 - INS GTGTACTGAAGATACAACAATGGCAACCAAAGGCAACTTAAAAAGGCAAACGAAGTACTTTTCAACAATAGCTTACACTGAAACTCGCGGAGAGGCGACGCTGCGCGCGAATTATCAGTAAAAATCTCGTAACAACCCATCTGCCACTTTTAGAAGGAATGGAAATTCTCAAAAAATGACGGAAAATAATAGAACAGGGTTCCTAAACGATGCATTTCTAACAAGTAGGATAGTCCAAAAGGGAGGATGCAAATTCTTTGTTTTCCACGCAGTAAGATATGATCCCAAGCTTTCGAATATAAAAAGGGAAGGATCGCTAGGACAGATCAGTTTTTAGCCCGTTTACTTATCTCGTTCCCTACTCTTGTTCTGATAGAAACCAGCAACAAAAACCTATTCACTCGCTTATTAATACCATAAAAAATATGGCTTACTCTAAAATCACATTACTAGCCGCTCTTGCTGCTATTGCTTACGCT tpg|BK006948.2|:342861-345467 7X4=5I17= 240=7X 
 tpg|BK006948.2| 383613 + tpg|BK006948.2| 383775 - INS CCTAAACGCGGTCTAAGCTCTGAAAGAGAAACGGAAACTCGACGTCTTTCCTCTGAAGGAAGGTTAGTCGTGGCACTATTTTTTCGCGTAGCTGGGGTACTATTTGAGGGAAAATATGAAGCTGCCGGTTGGCTAGTAAATGTAGATGCAGTAGTGTAGGAAGATTCAAATGGTGCGTGTGATGCAGTGGTGTATGGATTAGAATTGAAGTGACAGTTTAAATGAGTATCTGATAGTTGCGGTCTAAGCTGGTATGTGTTCAGT tpg|BK006948.2|:383071-384317 7X4=140S 69=1X178=7X 
 tpg|BK006948.2| 501544 + tpg|BK006948.2| 501873 - INS CCTCTCCGCTTTCATAATTATAAACGGCATCCTTCACTGAACCGTTTTCATCACTGGAACCTGGCAATGACGATTGCAAAGAAGCTGTATATCTCTTGCTCCGCCTTCTGGGAGTATTGTTCGCAGAAGTCGAGTTTATAGTTGTGACACGATAGATAGAATGACGTCTGTCAATTGAATTAGGTAACGAC tpg|BK006948.2|:501148-502269 7X159= 168=7X 
 tpg|BK006948.2| 63702 + tpg|BK006948.2| 63875 - INS GCACTGTTGGTTTCTGATAGGAGAACATGTTTTGGAATGTACTTTCTTGCCAAGGAATAGATGCGAACTTCAGCTTCGTCACCCATTGACGAGATTCCTAGTAATGAATTATATATATTACTACTATAAGCAGGCTTGAACTTCAATTTAGTGACTGGATAGCCCGTATTAATTGTTAGTTTGGGAAATGCCAGCGAGCCGCTATTGTTCAAGGACGTATTGGGGGCATGTAACGAGGGAGAGTTCCCGTAATTGAGGACTGTATTTTCGGCGGCATTGGCATTGTCGCCAACAAACCAGAGGCAGCATTTACCGTCTCTACCACCTG tpg|BK006948.2|:63032-64545 7X157= 72=1X235=7X 
 tpg|BK006948.2| 332779 + tpg|BK006948.2| 333230 - INS TATTAAAGGTATAGAGTATGTTACTAAGGAGCATATAGAATCGTCGAAGAAAAAGAATAAAGAATTCAAAGGATCGACTGCCAATCTTTCTTTGGGAAGTAGCAAATCGCTAGCTATGGAAATGGCTGTAAATGCAGCTGTAGATAGCGGTGTCCATT tpg|BK006948.2|:332449-333560 7X5=74S 68S11=7X 
 tpg|BK006948.2| 129415 + tpg|BK006948.2| 129719 - INS ATATATGCCTAGAATAAGGTATGAAACATGACAGATGGTTAACGATCGACTCGACACATTGTTGATGGAATAATTGGTCCCTAGTTAAACAGCGGAGAAATAGCCGCCCAGGATAATCGGAGAAAAGTCACGTGCAAAAAGAAATCATATTCGACGAAATAAACTAGAATAACTTTTGACGTTTAGCAATAATAACCCCAAATGGAAGCGAACATTTCCCGATCCTTTTAG tpg|BK006948.2|:128939-130195 7X6=109S 109S7=7X 
 tpg|BK006948.2| 385428 + tpg|BK006948.2| 385165 - INS AATCATTCCAATTCAGTTTGATAGTACCTTTTTTTTAAAATTTTTGAAAGAGCTATCGCTTAGCTATCGGCGGGCATATTGAATTGCGCAGTAGATGAAC tpg|BK006948.2|:384951-385642 7X25=25S 1S1=60S 
 tpg|BK006948.2| 527593 + tpg|BK006948.2| 528258 - INS GACTATCTATCGTTGTCATCTGTGACTAAAAATATACAGGAAAATAAACCATTGGCGCAAAATAGACGAATTCCACCACCAGGTTTTAGTCAAAATATATTAACTCCAAAAAGTACCAGTAACTTGGCTTCGCCTATGTCTTCTAAGGTTGATTTATATAA tpg|BK006948.2|:527257-528594 7X8=102S 141=7X 
 tpg|BK006948.2| 133193 + tpg|BK006948.2| 132533 - INS AGTGATTATTCCAATTTAGCTGGATGACAGCTCACAAAGGCAACGCTTTTATTGGAATCAAACATGTTGACAAAATATTTCTGCATGGCATTTTTCAGATCTGTTTTGGTAACATTCTGCAACCTTTCCAAATACAATTCATTGAAGTTGTTCCCCCTTTGCAAACAGAATTCATCAACATATTTGGACAGGGCTGTTTCAAAG tpg|BK006948.2|:132111-133615 14S95= 102=7X 
 tpg|BK006948.2| 648859 + tpg|BK006948.2| 649365 - INS CCTTCTGATTCACTTTACAAATTGATTAAGGAGACTCCTTCGGACTATCAATGGAACAAATCTACTAGAGCGCTAGTACACAACCTGGCATCTTTTGTCAAAGGTACAGATCTACCCAAGTCTGAATTAATTGTTAACGGCATCATTAATGGTGATTTGAAGACATCTCTGCAAGTCGATGCCGCATTTAAATATGTAAAGGCTAATGGCGAGGCATCCACCAA tpg|BK006948.2|:648397-649827 7X11=1S 112=7X 
 tpg|BK006948.2| 52187 + tpg|BK006948.2| 52640 - INS GTATACCGTAATATTATCTTTTCCTATAAAATGAATAATTTTTCATTCAAAAAAAGTTCGATTACGGGTAACGAGCAAATAGTTACTGTGAAAATTTTTAAGAATTGAGCGATGAGCTAAAATGTCAATGTCAGTCAATTAACAAAGTATACAATAGGCCCATATCATTTTAGATTGTACCTGAAGTGAGAACTAGGTAATATACGACGATGGATAGTGTAATTCAAAAAAGAATTTTTG tpg|BK006948.2|:51693-53134 10S117= 120=6X1S 
 tpg|BK006948.2| 252607 + tpg|BK006948.2| 253244 - INS ACAACCCCCATTTCTGGTCTGATTTCAACTTGGTTGAAAGCCTTACCGTTGTAGATACCGACGACGGAACCGATCATTTCTGGAACAATGATCATGTTTCTCATGTGGGTTCTGACT tpg|BK006948.2|:252359-253492 7X9= 103=7X 
 tpg|BK006948.2| 548300 + tpg|BK006948.2| 548593 - INS TGCTTGCGCAATTTTTTTAAATCCTTGTCCTCATGTTTCTTCCCCTTTAAAACTTTTGGTTCATCATCGTCATAGTACTCGCCCTCCTCCTCGTCATCTTCTTCAGATCCGCTTGAGCCGTCTTCTTCATCATCTGAGAATTCCTCTGTGCCAGAACTACATTCGTGGTCAGCGTTATCA tpg|BK006948.2|:547926-548967 7X82=53S 2S1=12S 
 tpg|BK006948.2| 365880 + tpg|BK006948.2| 365918 - INS GTCATTAATGCTGGATTGAATAGTCATTCACTGACACCAAGCTTTGCACATTTATCTAGGCGTAACTCATATAGTCGCCAAACATCTTCTACATCGCTGAAGAACGATTTGGAACTGACAGATTTAAGCAGAGTTCCCTCGTATGATAAAGC tpg|BK006948.2|:365562-366236 8X24=1X60=28S 34S4=7X 
 tpg|BK006948.2| 839866 + tpg|BK006948.2| 839599 - INS GTATATATCTATTAACCTGATCTCTGATCCAATCAAATTTTTATCGATGCTTTGAAATAGTTCATTTGTTTGTTTGTCAATCGCACTACCTTCATCAAGGTATCCTCTCAGCTTTTTTAGTTTTTCATAATATGCTGTGTTAGTAGTTGAAG tpg|BK006948.2|:839281-840184 7X3=174S 3S140=7X 
 tpg|BK006948.2| 735828 + tpg|BK006948.2| 735407 - INS GTCATATTCTCAGAGTCTCGCAAGTCAAGAAAACAGCTCCACAAAATGATAATATCAGTCAAGATTGTGACCTTCCGCATAATGGTGACCTTACTTCCATTACCATGGCTGTATCCGAGCCGTTTATTGTTTACCAATTACAATACAAGAATTGGTTAGATTCATGCGGCGTAGATATGAATGACAT tpg|BK006948.2|:735019-736216 7X8=4S 94=7X 
 tpg|BK006948.2| 564597 + tpg|BK006948.2| 564820 - INS ACTTGAATCAATAAACTTATATAT tpg|BK006948.2|:564535-564882 7X10=2S 8S4=7X 
 tpg|BK006948.2| 624945 + tpg|BK006948.2| 624254 - INS TTCATGCATCCTTGGAT tpg|BK006948.2|:624206-624993 7X1= 11S5=7X 
 tpg|BK006948.2| 155250 + tpg|BK006948.2| 155350 - INS TAAAGTGTT tpg|BK006948.2|:155218-155382 7X4= 1S4=7X 
 tpg|BK006943.2| 526927 + tpg|BK006943.2| 526735 - INS GGTGTACAATTTTTTACTCTTCGAAGACAGAAAATTTGCTGACATTGGTAATACAGTCAAATTGCAGTACTCTGCGGGGGGTGTATACAGAATAGCAGAATGGGCAGACATTACGAATGCACACGGTGTGGTGGGCCCAGGTATTGTTAGCGGTTTGAAGCAGGCGGCGGAAGAAGTAACAAAGGAACCTAGAGGCCTTTTGATGTTAGCAGAATTGTCATGCAAGGGCTCCCTAGCTACTGGAGAATATACTAAGGGTACTGTTGACATTGCGAAGAGCGACAAAGATTTTGTTATCGGCTTTATTGCTCAAAGAGACATGGGTGGAAGAGATGAAGGTTACGATTGGTTGATTATGACACCCGGTGTGGGTTTAGATGACAAGGGAGACGCATTGGGTCAACAGTATAGAACCGTGGATGATGTGGTCTCTACAGGATCTGACATTATTATTGTTGGAAGAGGACTATTTGCAAAGGGAAGGGATGCTAAGGTAGAGGGTGAACGTTACAGAAAAGCAGGCTGGGAAGCATATTTGAGAAGATGCGGCCAGCAAAACTAACTCGAGTAAGCTTGGTACCGCGGCTAGCTAAGATCCGCTCTAACCGAAAAGGAAGGAGTTAGACAACCTGAAGTCTAGGTCCCTATTTATTTTTTTATAGTTATGTTAGTATTAAGAACGTTATTTATATTTCAAATTTTTCTTTTTTTTCTGTACAGACGCGTGTACGCATGTAACATTATACTGAAAACCTTGCTTGAGAAGGTTTTGGGACGCTCGAAGTCTTCCGCTTCCTCGCTCACTGACTCGCTGCGCTCGGTCGTTCGGCTGCGGCGAGCGGTATCAGCTCACTCAAAGGCGGTAATACGGTTATCCACAGAATCAGGGGATAACGCAGGAAAGAACATGTGAGCAAAAGGCCAGCAAAAGGCCAGGAACCGTAAAAAGGCCGCGTTGCTGGCGTTTTTCCATAGGCTCCGCCCCCCTGACGAGCATCACAAAAATCGACGCTCAAGTCAGAGGTGGCGAAACCCGACAGGACTATAAAGATACCAGGCGTTTCCCCCTGGAAGCTCCCTCGTGCGCTCTCCTGTTCCGACCCTGCCGCTTACCGGATACCTGTCCGCCTTTCTCCCTTCGGGAAGCGTGGCGCTTTCTCATAGCTCACGCTGTAGGTATCTCAGTTCGGTGTAGGTCGTTCGCTCCAAGCTGGGCTGTGTGCACGAACCCCCCGTTCAGCCCGACCGCTGCGCCTTATCCGGTAACTATCGTCTTGAGTCCAACCCGGTAAGACACGACTTATCGCCACTGGCAGCAGCCACTGGTAACAGGATTAGCAGAGCGAGGTATGTAGGCGGTGCTACAGAGTTCTTGAAGTGGTGGCCTAACTAC tpg|BK006943.2|:523935-529727 601S64=2D38= 23=1X64=616S 
 tpg|BK006943.2| 745751 + tpg|BK006943.2| 745527 - INS ATACTGTAGCATCCGTGTGCATATGCCATATCAGTATACAAGTGCAAGTGAGTATGGCATGTGGTGGTGGGATTAGAGTGGTAGGGTAAGTATATGTGTATTATTTACGATTATTTGTTAACGTTTCAATATGGAGGGTAGAACAACAGTACAGTGAGTAGGACATGGTGGATGGTAGGGTAATAGTAGGGTAATGGTAGTGGAGTTGGATATGGGTAATTGGAGGGTAACGGTTATGGTGGACGGTGGATGGTAGTAGTAAGTAGAGAGATGGATGGTGGTTGGGAGTGGTATAATGAAATGGGACAGGGTAACGAGTGGGGAGGTAGGGTAATGGAGGGTACGTTAAGAGACAGGTTTATCAGGGTTGGATTAGAATAGGGTTAGGGTAGTGTTAGGGTAGTGTTAGGGTAGTGTGGTGTGGTGTGTGGGTGTGGGTGTGGGTGTGTGTGTGGGTGTGGTGTGTGGGTGTGGTGTGTGTGGGTGTGGGTGTGGTGTGTGTGTGGGTGTGTGGGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGGGTGTGTGGGTGTGGTGTGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGGTGTGGGTG tpg|BK006943.2|:744099-745750 7X475=8I26=21S 1=401S 
 tpg|BK006943.2| 47713 + tpg|BK006943.2| 47772 - INS GTATGGTGATGGCTGGAGTATGGTGATGCTGCTGTCCATGATGTAATTCTCCTTGGCACTTCGTAAAATTATTATTTGTCTGCAACTGGGGCACTAAAGCTCCACTACTTTCTTGCCGTTGCAATTTAACTATATTCAAAAGTTGTTCAGATAATACAGAGGTCTTCTCGTTAAACTCTTTGAACAATTGGTTCAATACTTCAAAAGTACGTTTACTCGCATTTGAAGCACCCTTCAAAAGTGATAATATTTCACTGCCAAGCTGCGTAGCGT tpg|BK006943.2|:47153-48332 104S113=4S 3S253=7X 
 tpg|BK006943.2| 659834 + tpg|BK006943.2| 660593 - INS GAATATTAGGTATGATGAGGACTCAATGTGATAACTGTCCATATTAGGTATGATAGAAGGAAGATGAATAAATGAAAAAAATGGATGGAATTCTTCCTTATAGTAAGTCACATAATCGTTCAATTGACTAGTTGTGGGGAAGGCTCCTGAATCGATATTATTGTCGGCTAGCATCATACTCCTTAGCTCATTGGTAAAAAGCACTTGAGATACTGAAGGGACAGAAAACGGAGATAACAAATCCGAAGGAGTAAGAACAGGCAGCTGTTTCTGTGTTGCATTAGAATCAGTTTCGCCGGGGAAAGACAAAGTGAGAACATCGTCGTTCACATGAGAATTATTTTGCTCTGTCCCGTTTAATACCTTGGAAATATCCAATTGCCTTGAGCTGAAAAAATTGGATAGATCGTAGTCCATCATGACGCTATCACGACGCCTCTTATGAGAACTATGGGAA tpg|BK006943.2|:658906-661521 7X161= 1S428=7X 
 tpg|BK006943.2| 548425 + tpg|BK006943.2| 548642 - INS AGATCAAGGCTTGTTGTCACAAGAGAGCAATGACGGAAATATTGACTCTGCTCTGTTGAGCGAAGGGGCTACGCTAAAAGGGACTCAAAGTCAGTATGAAAGCGGACTGACGTCTAACAAAGATGAGAAAGGAAGTGATGACGAAGATGCGTCAGTGGCTGAGGCTGCTGTTGCCGCTACCGTCAATTATAC tpg|BK006943.2|:548027-549040 7X166=14S 1=212S 
 tpg|BK006943.2| 551179 + tpg|BK006943.2| 551548 - INS GTACTGGACAGACATCATAGAGACAGGCGATTTTTCTCAATCGGACATAATCTCCTAAATGACCCTCAGGAGTTTGAGGCAAGATTGAATTCTTTGATCAGAAATTTTCAGAAATTTGTTAAGGCTAACGGATTAATTTCCTGGCTATCGCATGGTACATTGTATGGATATCTATATGATGGTCTGAAGTTTCCCTGGGATGTCGACCATGATTTACAGATGCCCATTAAACATTTACATTACTTGAGTCAATATTTCAACCAATCCCTAATATTAGAAGATCCAAGAG tpg|BK006943.2|:550587-552140 28S264=5S 59=1X211=7X 
 tpg|BK006943.2| 110538 + tpg|BK006943.2| 110540 - INS GGATATGGGATTTCCTTAACAAAGAAAACAATTCTCCACCTTCAATATAATCCATAATCATGAAAATTTGCTGAGCATCTTGGAAAGTCCCCCACATTCTAATAATAAACGGATGTGTTACGATAGAAAGCATCAATCGCTCGTCGTTGGTATGCTCCACCTGTTTCAATCTTACCACGATTTCCTTTTTCAAAACTTTCATGGCGTAGTATCTGCCATTATGTCTTGATCTAATCAAATGGACCCTACCAAAAGAACCCGTACCCAGTGTCCTTAATATCTGAAAGTCTTGTAAACTATACTTCCCACTTGTAACTCTCGCTTGGGC tpg|BK006943.2|:109868-111210 7X191= 164=7X 
 tpg|BK006943.2| 407736 + tpg|BK006943.2| 407826 - INS ATTATTATCCCGTGACGGGACTACAACAGTTATTATTCTAGCTGGTGAGATTTTAGCTCAGTGTGCACCTTATTTGATTGAAAAAAATATTCACCCTGTTATTATTATCCAAGCCTTGAAGAAAGCACTGACTGATGCACTAGAAGTTATCAAACAAGTAAGTAAACCTGTCGATGTGGAAAATGATGCCGCTATGAAAAAATTGATTCAAGCCTCTATCGGTACTAAATATGTCATACATTGGTCAGAGAAAATGTGTGAATTAGCTCTAGACGCTGTTAAGACTGTCCGTAAAGACCTGGGACAAAC tpg|BK006943.2|:407104-408458 7X5=159S 290=7X 
 tpg|BK006943.2| 36192 + tpg|BK006943.2| 36668 - INS ATCGCTCATAACGAGGAGAGATTGCCGAGATAACTGAGAAGACGTAATCTAAAGGCAACGCAGCATGTCTCGAGTTGCACAGCTCGACTCGATAGCGCTTGATAAAGAATTGTATGGACAGTTTTGGTCCGAGTTCAATGCAGCATTCAATACGAGTGAACACAAAGAGGAATGGGAGTTGGCACTGAACACAGTTGTGTTTATGTGCGCGACGAGGTTCCTGCCACACTATGGCTCTAGCTGTACGTATGGATC tpg|BK006943.2|:35668-37192 7X200= 128=7X 
 tpg|BK006943.2| 101304 + tpg|BK006943.2| 101330 - INS GAACCCTTGCAGCGACACTCGTCCTCGACTTGTTCCGTGTTCACGTTTAGGAAAGACGACGGCATACCGTCTTTGCTCTCGTAATATTCTTCGCTGTTGCTATCACTGAAATTCTGCATGACGCGAATCTCTTGGAGGACTTCTTCCTTTATGGGTAGCACCGTTCTTTTAGTTATGGCTTCATATTCATAAAATCCTGGGTATTCGTCTTCTTGCAAGTCGTGGAATTCCAATTCATGTGGTTGCCAATACTGTAAGAACCACCAGGCTAAAAG tpg|BK006943.2|:100740-101894 7X79=1X181= 140=1X117=7X 
 tpg|BK006943.2| 25361 + tpg|BK006943.2| 25399 - INS TTATGAGGTGGTTGATAACCAGGTCAACAATAACCTTGATACCTCTCTTATGAGCTTCTTCTATCATTTGGAAACAATCCTCATTGGTACCGTAACGTGGCCAAACCTTCTCATAGTTGGCAATATCGTAACCCATATCTTCTTGAGGAGAGTCATAAAATGGGCACACCCATATCGCATCGACACCTAA tpg|BK006943.2|:24967-25793 14S28=60S 92S3=7X 
 tpg|BK006943.2| 192002 + tpg|BK006943.2| 192746 - INS CCTCTCAAATATGTTCTACCCGCTGACTCGTATTTCAAGTCGAAGATCAACCAACTTGTTGGTTCTAAAGGTGAGAAAGTTTTCGGCATCAATTTGAATGATTTGGTGGCAAGACATGAAACAAAGGATCCAGTGGTGAACAATACGCATATCATCGTTTATAGAGAAACGCCCATTGCATTGATTTCGTTAGCCCCTAACATGACATTAAGTACTGATGAAAATTTAGTCATGAGTGTTACTACTG tpg|BK006943.2|:191494-193254 7X278= 7S225=7X 
 tpg|BK006943.2| 484612 + tpg|BK006943.2| 484666 - INS TTCCTATATCCTCGAGGAGAACTTCTAGTATATTCTGTATACCTAATATTATAGCCTTTATCAACAATGGAATCCCAACAATTATCTCAACATTCACATATTTCTCAGTTGCCTTACTTTAACAGAAGATAACAGAAGTGAAGAACTTATATATTCTGATGAGTCTTTCATATTAGCCAATTCTGAATTTTCAGTAGATGATCTAGT tpg|BK006943.2|:484184-485094 7X4=99S 95S7=1X1=7X 
 tpg|BK006943.2| 113293 + tpg|BK006943.2| 113706 - INS GGCGTACTTACCTGATGTTAGTAAGATAACATTCGATTATTTCAGTAGTTTATTGAATTTCCATAACTAAATATATATTTAAGATATTAATAATTGAGACATGAAATGTACTGACTAGATACTTTTATATATTTTACATTATTCATTCAAATTATTTCCATCCTGGCGTAAGGACGACGGGTATATGCTCATTAAGAAGAGCGTTCGATTATACTTTACCGTCACATCTTTCGGAAAAAATTTTAATGACCTGCATCTGTCTTTCTTGTAAGATGTTCAATTTGTCCATTAAACTTTTATCAAATTCTAGGTATGTTTTCCAAACCATAATACTTTGCTTTTGGGTTAACATATCACTGAACTGCGTATCTGCTCTCAGGCGCTGTAATGATACTTGATGTATTGTTTCTTTAAGTTTGTTACATTGGTTATTAAACAGCTGCACGTTAAGC tpg|BK006943.2|:112375-114624 7X216=2S 12S416=7X 
 tpg|BK006943.2| 641388 + tpg|BK006943.2| 641893 - INS GCACTACACCACGATCCGTGACCCACTGCTGAAAATTGATTTCAATGTCCACACCGTCTCGATGATCCAGGCTGTCGTCTCGAACACCGTCCTGTTGCCCACCCTCACGACGCCAATGCATTATAATGTTGTCACCTACACAGATTCGTACAGTTCAATGGTATCTTCCCTCAGCGCAGGGTACTTT tpg|BK006943.2|:641000-642281 7X4=306S 94=7X 
 tpg|BK006943.2| 123219 + tpg|BK006943.2| 123393 - INS GGGCTTGACTATCGGTGGCTTGAGCAGTAGCAGCAGAAGTGGCTTGGACTTGACCGTCACCAATTTGAGAGATAACGTCTCTCTTAGCTTTTGAAGAGGTAATAGCTTGAACAGCAATACCAAAGGTGGTAGTGTATTCGGCAGCACCACAAGAGATGGAGCCGGTTGGGGTTAAGGTGGACCATGGTTCACCTGGAGTGTAACCTTCAGCAGAAGCAGTGGCGGATAGAGCAGCAACGGAGGCAGCTAGGGCGACGTTTTT tpg|BK006943.2|:122681-123931 7X3=196S 131=7X 
 tpg|BK006943.2| 108890 + tpg|BK006943.2| 109131 - INS GATAGAGTCTGAGTGATTTCTTCCCCTCATGTATATTCTATTTCCTGTACCATTACCAACATTGTTGGTGGCATTTGAATTCATTCCACCATTTCCATTTTTCATTGGTGGTGACCTTGGTGTGGACAAACTGTTCTTCCTACTTCTTGTGCGATTGCTATGATTACGTACGCCCAGACTGTTTCTCCTTCTAAGTTTTGATTCTTCGTCATAATCAAGCATAGCATCAATAGAAAAGTTATTTTCCTGATCCAAAACATGGTTGGCTGCAACATCATTGCCGTTCTCAGATATGTCTTTCTTTGTCGGTTGATCAGATTCACCTTGTTTTATATTAGCCTCACTTTTGGGATGAGTTTCGTCACAAC tpg|BK006943.2|:108140-109881 7X267=55S 187=7X 
 tpg|BK006943.2| 138347 + tpg|BK006943.2| 138386 - INS GGATAAGGATCAACTGGGATTTGGACTCTACCTTGCAAAGGTCCATTCTCAGCATCCTTTGCAATCAGGGCAAGTCCTTGCAAAGACTAGAAAACGTCACTGACCCGGCTTGTAACGATATCATCTCCAATGGTCACTTTTCCAGGAGCAACGTCT tpg|BK006943.2|:138021-138712 7X4=74S 74S4=7X 
 tpg|BK006943.2| 31237 + tpg|BK006943.2| 30520 - INS GTTAAAGACCTCTTATTCAAATTTTGAGGGTCGGGAGAATTAACTCGTTAATTATTCCTGGTGTCGAATTTGCGTCATTCCTAAACTTGGATATTCTTATATGGCAAAAAAAGAATTTTTTATGCCACCAACACGACGGCATATTCTGGAGTGATTATAGCCACTGCTAACAAGATAAGGCGGTAACACCCGATTGTGCAGATGTCCTCATTTATCCTGTTTCCGAGCATTTGATTAACCGTCTCTGTGAGACCAGTTAAAGACCTCTCTCAAGAAAAATATGTAAATTTTTTTCAGCCACTTTATCGGCACTGGAACGAAACGATATGGTATTCCCAGTATCAGCCACGGCCCCGTGTAAGCCGTAAAGTAAACAAAAATTTTTACCACTAATTTCGTTGCGTATCAATTTATACTATTCTTTGTGAAAACCTACAC tpg|BK006943.2|:29630-32127 7X5=186S 411=7X 
 tpg|BK006943.2| 500709 + tpg|BK006943.2| 500731 - INS TATTGCATTCTGCGAAGACCCTTTTAAAACCTGAAACAAATTTATTGTATTGTGGCTCAATGGACTTTTCCAGATAAAATTCTACCCATTTCATGACAAACTCATGCTTGTTACTTTGGGTTATTGGCACATTTCTGCCATTTTCACATAATTCTACCGTTACATACTCTTTGCTCGATTTACTGTCATTTAAAATCCAGTTGTTATTTCGATACGTAGTCTCAAATGTTAAAGAAAAGACGTCTTCGAAATTATCCTCTGTGT tpg|BK006943.2|:500167-501273 8X156=41S 2S1=185S 
 tpg|BK006943.2| 42558 + tpg|BK006943.2| 42561 - INS CGCCTGTATACCCAAATATCTCTACGAAATTTAACCAGACCGGTTCATATAACTCAATTTTCGTACTTCTTGGTTCAATGAGACTATTTTCTTTCGAGTCATTCTTTACTTGCACAGTAGAATCATTATCGTTATACTTTATCATCATGTATTCACGTAAAGAAATGATCCATAATGGGACTAAAA tpg|BK006943.2|:42172-42947 7X196= 8S167=7X 
 tpg|BK006943.2| 699555 + tpg|BK006943.2| 699768 - INS ATCAAGATGGCATCCAGTAAAATCAGCCTAGTTTCTGTAACATGCGCAGTATCGATTGCAACCAAGAGAGATGCAAACGCACATGTAATAGCCCTGAAATTCAGTTCCTTCAAAGTGTTGAACATAATTGGTACAGTCAATGTGCCCAATATCGCGTTGAAAGAACGGTACGCGATATATGGAGCTGGATGAGTT tpg|BK006943.2|:699151-700172 7X148=22S 4S1=347S 
 tpg|BK006943.2| 558820 + tpg|BK006943.2| 559208 - INS GCCCGGTTCTTAAACTACTCCTTGGAACATGAATTGTCGATAGAAGAGTTCCAAGCAGTTTCAAATGACATAAACAATAAGATTTTGGAGCTGGTCCATACAAAAAAAACGAGCACTAGGGTAGGGGCTGTTCTATCCATAGACACTTTGATTTCATTCTACGCATATACTGAAAGGTTGCCTAACGAAACTTCACGACTGGCTGGTTACCTTCGAGGGCTAATAC tpg|BK006943.2|:558354-559674 7X7=106S 108S5=7X 
 tpg|BK006943.2| 213439 + tpg|BK006943.2| 213861 - INS AAGTTATACATGTACTTGATCTGTTTCCTCGGTTATTTTATTGATAAACTCAAAGGTATTGTTCATAAATGTCAAAAATTCACTTTCCGAAAAATTCAAGACACCATTTGAAAACAAGACACGGGATTCTAGTGATTTCTTCTTTTCCGAGGAGCTCTTTGATGATGTCAACAATTTGATGATATCGAGTAAGTCATTCAAACCTGATAATTCCTCATTGACATGTAGATCAACGAGTAGGGCCTTAATAAACTCAATTAATATTCTTGCCTCGCCAATTTTAAAGTTGACTAAAGCTGAAGAATACTGTTGTGCAATCAAGAAAAGGAACGAGCCCAGTGCCTTTACTGGATCAAGTGTTTTGATTAACGTAGAAAATAATTTAACCCTCCTATGTCTTGGAACATGTTGCAAAGCGGTTGTGAAG tpg|BK006943.2|:212571-214729 7X170= 401=7X 
 tpg|BK006943.2| 591059 + tpg|BK006943.2| 590462 - INS CAATCATTTGCATTGTCATCATTACCATTGTTAGTTTCATTGTTACTTGTATCGTTTGCCCCAGCATCCGATACAATATTCACTATGTTGTTGGCGTTCCGGTTGGCGTCATTGTCATTATTGTTATTCCATGCTGATCTTTGGTGGGCTATTAATAGTTCTCTTTGTC tpg|BK006943.2|:590110-591411 7X95= 159=7X 
 tpg|BK006943.2| 219016 + tpg|BK006943.2| 218954 - INS GCTTGAGCTTGAAACAATCATACACTTTTCACTTGAGATGGAGGGGGTACGTATGTGGAGGTTTCAATAAACCCTTCGTTATCGTCGGATGAATTGTTTTCTGCATAATCATCAAAATGATCCACTGCAGGAGCCAGAAATGAATTTTTTGAACTTGAGCCTAACGTTTCGCCATCCGACGTACAATTTACG tpg|BK006943.2|:218556-219414 7X1=1X10= 10S170=7S 
 tpg|BK006943.2| 152030 + tpg|BK006943.2| 152641 - INS TTGGTATTGATGTATGTTAAATCTGTCCTCTAATGATCTCATTGAATCCAATGCCCCTTCTAATTCTGAATTTCTCACCAGCATTAAAATTGTTGCATTTTCTCGTAGGTGAAAAGAATCAGAATCATTCTGTCTGGTATAATTTAAAGTGTAGTCGTCGTAGCTATTGCGGGAAAGTTTTACTTTAGGAAAATAGTTTCTTCTTCGACTTGTATCATATTGTTCTTTTACTCTTTGGGAAAGAGCAGTATACGTACTGTCAATCTTTTGGTATTTTCGTATGAGGAATAACTCTTTGCCAAAAATATAGATCATAAAGGTCCATATTGGTAAGAATATGCCAACGATGTATAGC tpg|BK006943.2|:151306-153365 7X349= 333=7X 
 tpg|BK006943.2| 103559 + tpg|BK006943.2| 103537 - INS CCACTGCTGTCGTCTGGCCAACGAACCCTTTATTGTGGCGTCAATGAATTCTCCGTTCTGTAACATCATAAAATAAAAATGCTTGAAATGACGTTGGTCATAGTCTATTAACCTATCTCTAAATTCCATCTCCTCGATCACCTCACCTTTGTACTCGTAAATGAACTGGTTGGCTTCTATGTCCTGTTCGGCTCTTACGCCATAACC tpg|BK006943.2|:103109-103987 19S91= 53=58S 
 tpg|BK006943.2| 616003 + tpg|BK006943.2| 616167 - INS AAGGCCATTGTATGCTATGCTAGGATTGGGCCCTAATTGGGAATAATAATTGTTTTATTACTGCGTAGTCAAATATGTATTTACAGAATTCTTTTAAATATATAATTCACCTACTCATCATAGCCACCGCCAAAAGAAAGGAAACCTCCAGTTTGTCTGGAATGTCTCGAAAAATAATCGAAATCGATGGACACAGCGTTTGCTAATAACACGGCCCTTTGATCCAAAGTTAGTACTTGAGAACTTAGCATCTCAGTAGGATAAATATTATCAAAGCATCTCTGCGAATCAAATCTAACAACATAAACACCAGTATCGGTAAACATTTCTCTTCCTAAACC tpg|BK006943.2|:615307-616863 7X12=293S 320=7X 
 tpg|BK006943.2| 709778 + tpg|BK006943.2| 710147 - INS GCACGCGTATATGTGCTAAGGTTGCTGAGCTATTTTTTCTATACTATTGTCAAACTCCAAAGATATTTTGAGCTTTATTTTCTTGCAAACAAAATACCCTACTGCTTAATAAATGCAATGTATACATAGTTTTCAAGGTACATTATATTTTAAAGTTACCTCAGGCCTGTTTGCCCTTGCATTCTACAGTCCCTTTGTAAGGG tpg|BK006943.2|:709358-710567 165S43= 4S187=7X 
 tpg|BK006943.2| 248225 + tpg|BK006943.2| 248035 - INS CTACAGACCCTGATGAATGGACAATGCATCGCGTCACCTCATGGTTTAAATTTCATGATTTTCCAGAATCCTGGATATTGTTTTTCAAAAAGCATCAATTGTTTGGTCACAGATTTATAAAGTTGCTTGCATATGATAATTTCGCTGTTTATGAAAAGTATTTGCCGCAGACTAA tpg|BK006943.2|:247671-248589 7X5=354S 88=7X 
 tpg|BK006943.2| 252622 + tpg|BK006943.2| 253276 - INS GTGATCATCTCTAAATGGACATGATGAATAGAATGCACATCGTTGCCAACGGTGAAGGCTTGCTTCTGTCCAATTCATGGGTCCTTATGAGCACCCATCTTAATAGGTATTTTAAGGGAAAGAAATAAATCAAAAACCATGCAAACGTGATAAGCAGAATATAAACGGTATTGACAGGGCTCCCTTCTGCACTAGAAAGAATAATACTTAATGCTAACAAAATCCATCCCATTATATCGTTAATGATACCCGCCGCAAGGACAACGATACCTGCTCTATCCTTGAT tpg|BK006943.2|:252036-253862 19S5=1X125= 112=38S 
 tpg|BK006943.2| 608058 + tpg|BK006943.2| 608755 - INS AACCCGAGGGGAGACTAGAGAATCATCTCGGTTGAATGGAGCATTATTTTTTTAGTGGCGCCCGCCCGGAGAAATGGACGTTGGCGAATGAGCCATGAATTATTAACCGCCCATGTCTACCAGATACCACATCGTATGACAGTACCAGCCTAGTCCCGGTAAACCGCAAACGGACCTTAATTGTGACGAAGGGCCCAAATTTGATGGGTCGGTGTTAATGATTAGTCC tpg|BK006943.2|:607588-609225 7X56=1X42=15S 1S1=320S 
 tpg|BK006943.2| 665007 + tpg|BK006943.2| 665233 - INS CCTCAAGAACATTTAATTTTTTCTTGCCATCGTCTTGTCCTTGTACCGGTGCCAACTCTTGTAAGGGCTTATGAATAAGGAAATCACCCATGTATAAGGCAGCTTCCCATGTCCTGAAACCTGTAGTACTGGCCGCACTGATCAAATTCGGTGTTTCCTC tpg|BK006943.2|:664673-665567 7X5=75S 75S5=7X 
 tpg|BK006943.2| 121368 + tpg|BK006943.2| 122093 - INS AAGGGTCCTACGTCTATTAAAAAAAAAATATTTATCTAAATAAAAGAAACCTTCTTTTAGAGAACCTTAAAAATGTAATATACAAATCATTCATACCAAAATCTTTTTACAAATCATAATCTTTTTCTATTTCTTTTCCCTTATAAAAGGTAGAACATTAGTAC tpg|BK006943.2|:121026-122435 118S24=1X113=1S 82=7X 
 tpg|BK006943.2| 543782 + tpg|BK006943.2| 544551 - INS CAAAATACAGACCCGCATACCTCCTGTATATGAGTTTCGTCGAATCGGAAAACTCTACGAAGTTACTCTGATGCTTATGATCTCTGGAAGATATGAGTCTATAAATCTGCGCAATGGCATCCTGGCTACGCTGAGGATCCGAACTGTGTACATCGAACCATCTCACCAACCGCACCACACCCTGCTTATTAAAGCACAGTATAAACTG tpg|BK006943.2|:543352-544981 7X23=81S 8S1=189S 
 tpg|BK006943.2| 146524 + tpg|BK006943.2| 146623 - INS GTAGTATAGTATATGCATTTCATAACATGCCACTGTCAGTGGCGCCACGGAAGGATAGCGGGACTTTATCAAATCATTAATTTCTGTGCATAAAGTGTATAGTATATTCATATAGATATGTATATATATCATTGAATACAGAAATCTTCGGGTGTATACAAC tpg|BK006943.2|:146186-146961 7X210= 142=7X 
 tpg|BK006943.2| 448598 + tpg|BK006943.2| 448835 - INS CGGCTAGTAATATATATACGATTAATCAGACGCGTCTGATTAATTTCAAAAGTTAAAATATAAACTATTTTTGAAATCCCATTGCAATAAGCGAACTATAGCTGAATCTTTCCTGCAAAAATGGAAGTGAAGGGCAATGGACGCATTGTTAACAAAGTTCAACGAGGATAGAAG tpg|BK006943.2|:448236-449197 21S73= 45=49S 
 tpg|BK006943.2| 542679 + tpg|BK006943.2| 542971 - INS ACTTGGGAAGTATTAAGTCAGCATCATCATATGAAAATACTTCATAACTTTTCTGGAGGATACCTTTTGAAGAGAGAAACCTGTATTTTGCACAGTGGATTAGAGCCGAAACTTCATATGCTGCTGCGTTATTTTCCATAGCTATAGTAACGTTGGAACAAGAATCAACTATTACCTATCGAAGAGTTTTCATGTTACTATTATATTATCCCATACTGTGTAAGAAGATAACATAAGGATTGAGAAACAGTAACAAAGTCTAATGAAAGCTAAAAATGCAAGGATTGATAA tpg|BK006943.2|:542083-543567 9S269=1S 12S7=7X 
 tpg|BK006943.2| 297147 + tpg|BK006943.2| 296854 - INS AGAAAGATGATAATCATTAACTTTTAGAAAAGGAAATTTTGCCGACAATTCCACATAATGATCAGCCAATACTTGCATCATCTGATAAGTCTAATGGGACGTTGAAATCACTAGCTGGGAAAGTTAGTTCAAACAACAACGCTTCAAAGGAAGATGGCACTATCATTAACGGCACCATTGAGGACGATGGCAATGATAATGATGAAGTTGATACTACGGTTCGTATTGTTCCTCAAGATTCAGATTCCTCTAGTTTCCCAAAGTCAGATCTTTTCAAAATGATCGAAGGTGATGATACAGATCTACCGCAATGGTTTAAGGGCAAAAATTCGAGAACTTCCGGTAATTCCAAAAATTCAAAGCCTTACACAACGGTTTTGAATAAAGACATAGACAATTCTAAGCCAGATCCAAGAAATATTTTGCCCCAGCGAACCCCAATAAGTGCGGC tpg|BK006943.2|:295938-298063 7X4=156S 4S423=1X9=7X 
 tpg|BK006943.2| 28307 + tpg|BK006943.2| 28560 - INS TTTTTTTTTTTTTTGAGGAACCGATTAATTAATACATCGTAGCCTCTGCTTATTGCATAACACAACAAAAAAATACAATAATACGCAACTTTTGTTTATAGAAAAATAAAAATGGAACATATGATATTCTCTGTTCGTCATATGATAACTTAAGCACTTTCGTGTGTACATAGGTATTCTAGTGCATTGGAATGAGATCAATTATGATTTCCTAACCCAGAATTTATATTACTAATGATTTCAGAATTAATAAAAGCTGAAATAAAAGGAGTAGCAATGTAATAGGAAATAAACGAG tpg|BK006943.2|:27699-29168 7X222=37S 4S1=158S 
 tpg|BK006943.2| 366526 + tpg|BK006943.2| 366932 - INS CTTCAATACACCTCAACAAAACAAAACGCCCTTTTCGTTCGGGACTGCCAACAATAACTCTAACACCACCAATCAGAATTCCTCTACTGGTGCGGGCGCCTTCGGAACAGGTCAATCAACATTTGGTTTCAACAATTCTGCGCCAAATAACACGAACAATGCAAACTCTTCAATCACACCTGCATTT tpg|BK006943.2|:366138-367320 7X5=88S 88S6=7X 
 tpg|BK006943.2| 531156 + tpg|BK006943.2| 531877 - INS TTAAGAGAAGAAGGGATCAGTGCTGAAAATATCAAACAAAAATGGTACCAGCGACAGTCGAAGAAGCAAGAAGATGCAACAGACGAAAAAAAAGGTAAAGCGGAGGATGATAGCTTTACTGCCGAGATATCTCGAGTAGTTGAAGATGAAGAAATTGATGAAATTGGAACAGGTAGTGGT tpg|BK006943.2|:530782-532251 7X112=23S 1S1=184S 
 tpg|BK006943.2| 412407 + tpg|BK006943.2| 413031 - INS GAATTACCGGGTGCGTTTGTCATGGCAGCAACCAAAGCAGCGTCATCCTCATCATCCTCATCGAAGTCGTTATCTTCGTTATCGGATCTACCGGGTCTTGTTATTTCAATATTTGTTGGTAGTGGAGGTTTCCTGATATCAACATCCATTTGAGGTAACCAAAATGGGATTGAATCCACTTTATCATTTAGTAAGGTA tpg|BK006943.2|:411997-413441 7X5=94S 88S11=7X 
 tpg|BK006943.2| 462909 + tpg|BK006943.2| 463012 - INS TTTGCCATTAATATCAAGCCAAACGCCACGGAGACTCTATTTGAATCACTAATCAACGATACCGCACCACTATTCAATTCTACGCTGTTTAATCAGGTGGTATATGAAACTGGTAGAGACCCGACAAACCTAAAATCAACGATTTTACCGGTTGCTCAGACCATTGAAGAGTACTACCATACATTCTACACACTAAATTATCTGCCGCCGTTATTGACAAACATAACCCAGGTATATCGTTATGCACTAACTAACAATGCAAGGTATATCGC tpg|BK006943.2|:462351-463570 7X255= 209S7X 
 tpg|BK006943.2| 534587 + tpg|BK006943.2| 535334 - INS GGGTTAGGTAGACAAGAGCATTGGAAAAATTTTACCACGAGGAGAACAGGTGGTGTAAAAAGTTAGCCTCATGGTTTATACCCCGAGATGAGACCATTATCAGTGTTGATGAGGAAACAATCATGGATGAAAGTACGGTCAATAGCAAGAGAAAATCCTATATGTATGAAATCAGGAACATGGTAATCAATTCGACAAAAGATTAGCCCTTTAGCCTTCTTATAAC tpg|BK006943.2|:534121-535800 7X438= 212=7X 
 tpg|BK006943.2| 186762 + tpg|BK006943.2| 186974 - INS ATATTCTCTCCACGCAATCTTGAAGTATCAAATTTGCATATTGGTCAAAGGTTCTTAGTACACCGAATAGCATTCTTCCATCACGCAAAAGAACGAAGATTTTACGGTCTACTGAGCTTACAATAGCAGCGGTGGTAGTGAAGTTATACTGGTCGAGATATAAATCGGCCTCACCTTCTGAAA tpg|BK006943.2|:186382-187354 7X5=86S 88S4=7X 
 tpg|BK006943.2| 70658 + tpg|BK006943.2| 70748 - INS ATAGTTGTAACCGTTTGGCTGAGATGCAATGATATACGCAACATTGCATTCAAAGAAATTGCAAAAAAGACACAATAAAACGTAATTTGTACAAATATTTTACTATCATTAGCTACTGGATGCAGAATGGATGATTGTTAGGGGGAGGTGGGGTACAATTGTTTGTTTTTGATACATTTTCTCTTTCAAATCGCAACCAATTCACTCTGCTAATGTGATAACAATGGCGCCTGTCGGAAAGGTGAAAAAAAAAAAATGCAAACAAATAAATTGGCACGGTGTGACATAT tpg|BK006943.2|:70066-71340 7X272= 271=7X 
 tpg|BK006943.2| 433909 + tpg|BK006943.2| 434169 - INS AAATATAAGCGTTTGACACGTCTATTGTCCTCTTATAATCAACATTCTCCCAAGTCGCAGGTGGCTCGTATTGGGCAGCAGAAGACACGTTGAAAAAACATAGGAACAATCCCACAATCCAAGAGAACCAAACCTGCCTCATTTTTTCAGCACCAATATTTTGTAGTTTGCGTCTTGTTCCGAGCTAAAGAAGCAATCGGGTACTTGTCAAAGAAGTAGCTTGCTTAATAAAAAGCAAACATTAATTTGTTCTGCATACTTTGAACCTTTCAGAAAATAAAAAACATTACGCGCATACTTACCCTGCTCGCGAAGAAGAGTAACACTAACGC tpg|BK006943.2|:433231-434847 7X166= 199S3=7X 
 tpg|BK006943.2| 66795 + tpg|BK006943.2| 67160 - INS TATGGTGGGCACTATACCGCGTCTCTAAACTACAGGAAATAATCCAAAAGTCACGCCACGGATATGATGAGCGTATCAAAAAGATATACGATGAACAGATGAAGTTGTATGAATTTAATAAGACTGACGAGGAGGAAGATGTTTCTGATGATATGATAGAATGTAATGAAGATGTGCAGGCCCCTGAATATAGTAATCGTAGTTTGGAGGTTGGGCATATTGAAACTCAGGACTGCAA tpg|BK006943.2|:66305-67650 87S57= 209=7X 
 tpg|BK006943.2| 237094 + tpg|BK006943.2| 237736 - INS CCTATCCTATCACATTTGGACGCGAACTCGAGAGAATCCAAACTGGCTCAAGTGGGTCGTACTTTGTGTATGGAACACGGGCCGACGAAAGCGTTCCGGTGGGGGTCTTCAAGCCCAAGGATGAGGAACCATATGGCCCATTTTCTCCCAAATGGACCAAATGGGCACACCGCACGTTTTTCCCATGTCTGTTTGGCAGAAGTTGTCTGATTCCAAACCTCGGGTACATCTGTGAAAGTGCGGCTAGTTTGTTGGATAGGCGACTGGAAACGCATCTAGTACCCTATACAGATACTGCATCTATAGAGTCTTTTAATTTTTATGATAATAGAAAAAAATGGGTATTGGGATACAACCTTCAGAAGAAGAAACAAAAAAAGCTGGGTTCTTTCCAACTTTTTTTGAAGGAGTACATCAA tpg|BK006943.2|:236244-238586 7X309= 405=7X 
 tpg|BK006943.2| 619835 + tpg|BK006943.2| 619157 - INS GATCTTTGGATTTAAACAACCTTAATGGCAATTACTTTATCATTTTCATCTTTCAGCATTGTGGCCCTATTTCTATCGCATAGGGGCTTCAAACAATAATAGAGCAAGCTTTCGGGCATTCTATGGAACTCCCAATTGACTGTTTCATCACCTTCACTCAATTCGTATAACGTAAGGACTTGATTCAGTTTTCCAGAGTCTTCGAACCACTGTAGTATCAAAGAAGCCCAACTGTCTAAGCTCTTCCATAATATAAAATATCTCGTAG tpg|BK006943.2|:618607-620385 7X5=359S 159=1X92=7X 
 tpg|BK006943.2| 108005 + tpg|BK006943.2| 108529 - INS TTCACCTACAGACAAACTGTTCTTCCTACTTCTTGTGCGATTGCTATGATTACGTACGCCCAGACTGTTTCACCTTCTAAGTTTTGATTCTTCGTCATAATCAAGCATAGCATCAATAGAAAAGTTATTTTCCTGATCCAAAACATGGTTGGCATTACTATTTGCAGGGTTTGAAGAACCTGCGTTTTGTGGGAAGTTTTTCAGCCGTTCCCTTGGTTGTCTTTCAACCTCATCGCTACCAACTGTATAGCGG tpg|BK006943.2|:107485-109049 7X243= 56=1X181=7X 
 tpg|BK006943.2| 194533 + tpg|BK006943.2| 194535 - INS AGAGAGGTATCCATGACAGAGGCCCATCCACCAAATCCTAGCCAGTCCAAGGAAACTATACCGTTTACAGAAGGGAAGTCCGAACATTTGACAGTACCATCTTGGAATCCGCCATCACGCTTCTGTTCAGAGGTATCCTTCTCAGATGAGGACAATGTAGTGGTAGTAGCAGCAGATTCTACAGTACTAGTAGCGGCATTGGAATCTATGTATTGAGTGACAGTGACAACCGCTGGTTTTTCATCTTTGTGATGATCTTCATGGTGACTGTCCGCTGGAGCAGGTGCAGGGGCAGAAAATGCGACAGAAGAAAGGGAAGACAATATTAAAGCTGCGGAAATTTTCATTATGTGTTAGAGAGAGA tpg|BK006943.2|:193791-195277 7X6=177S 353=7X 
 tpg|BK006943.2| 342615 + tpg|BK006943.2| 343287 - INS CTAGAGCATAAGAGGAGGGATAAAGAAAGAGGTGTTGTGTGGGAAGAAACGATTATTTTACTGCCAGATAAGGTCCGTTACGTGTTTTTATCGGCCACCATTCCAAATGCAATGGAGTTTGCTGAATGGATATGCAAAATTCATTCTCAGCCATGTCATATTGTCTACACAAATTTCCGTCCAACTCCTTTACAACATTACCTGTTTCCAGCCCATGGAGATGGTATTTATCTGGTGGTTGACGAAAAAAGTACCTTCAGAGAGGAAAATTTCCAAAAAGCAATGGCGTCCATAAGTAACCAGATAGGTGATGATCCAAATTCCACTGATTCAAGAGGTAAAAAG tpg|BK006943.2|:341911-343991 7X199= 324=7X 
 tpg|BK006943.2| 322858 + tpg|BK006943.2| 323015 - INS TATGACAATCAAGATACCAAAATTCAGTCATGTTTAAAAGGGGAAGGTACGATAGAGATATATATAAAGTGTTCAATTTACTATAATTGCGTATAGAATCCATTGTTACTTGCTCTCAATGAAACAACGATTCATTCGTCAATTTACGAACCTAATGTC tpg|BK006943.2|:322526-323347 7X80=39S 4S1=171S 
 tpg|BK006943.2| 421178 + tpg|BK006943.2| 421809 - INS AATAACAATTTCGATGCTTACATTTTATGCTAGTATACACCACGCATATGTCTGTCAATGTACCTATTACAGAAGGAAATGTTCAAGAAGCAGTTCAGACAGTACCGAAGCAGAATTAAAAATCCATTATTTGAATATGATCTGATAGTCATATATATGAGCAATACAGGTCTTCACATTAAATGTATGAGAACTGCCGGAACCACTATTACATTGGTCACAATTAGGAATGAACCAATCGGCGTGTGTTTTATATCCCCCTTATATAAGTC tpg|BK006943.2|:420620-422367 7X194= 136=7X 
 tpg|BK006943.2| 189019 + tpg|BK006943.2| 189201 - INS GTGTAATTCCATTATTGTTAGGATGGCCCCATTCATCTACAAATATTCTGATTCCTCCCTCAACTTGTGAGCTTAGAACTTGATCAAACTTGCTTTCAATATTGTATTGTAATGAGGGATAGTTAACCAAATCATGGACTAGATGAATTCGCAGCACCTCTTCAGTCTCACCA tpg|BK006943.2|:188659-189561 7X4=6S 8S155=7X 
 tpg|BK006943.2| 725701 + tpg|BK006943.2| 726037 - INS CAATACAATATACGAATCATGGCAAGGCTCACCGTTTCCTAAGGAAACTACTGTGGCAACGAGATCGGTTTTACACTCATCTACAGTCTTAAAGGATGTGGTATGCGACCGTATGTTTTGTGATATCTCAAAACATTTTTTGAATGAAGAAAACTACTTTGCGGCGGGAAAGGTGATTAATAAATGCACTAGTGATATTCAACTGAACTCCGGTATAGTCTACAAGGTTGGCGCTGGTGCAAGTGACCAGGGCTACCAC tpg|BK006943.2|:725169-726569 7X6=152S 243=7X 
 tpg|BK006943.2| 700950 + tpg|BK006943.2| 701040 - INS ACTGCTACAGAAGTACGGTCTTATTTGCCATGGTCAATTGATCAGTGTGGCAAGAGGCGAACAAGACTATTTCAACGAAGCCGGCATACCAACTGCTACAGAAGGTTGCAAAAGTAATGCATTAATGAGGTGTTGCAAAGATCTCGGCGTCGGTTCTGAATTATGGG tpg|BK006943.2|:700602-701388 7X4=79S 80S4=7X 
 tpg|BK006943.2| 460247 + tpg|BK006943.2| 460901 - INS GTTTTATTTGTATCCCAATAGCAATTTTTATATACTACAATAAAAGAAACCAGGGTCCACGAACACAACTTACATCGCTACTCAATATCGGTTTGAGTACTCTAACAACTTTGCTTGGATGTGGTTGGGCAATGTACAAGATATACGGATACGAGTTTCTGGATCAGGCATACTTGTACCACTTATACAGAACGGATCACAGACACAATTTTTCAGTGTGGAACATGCTATTGTATTTAGATTCTGCAAATAAGGAAAATGGTGAGTCCAATCTCTCAAGGTACGCATTTGTGCCTCAATTGCTGCTTGTTTTAGTAACTGGATGTCTTGAATGGTGGAATCCCACATTCGATAACCTATTGAGGGTTTTATTTGTGCAGACGTTCGCATTTGTGACATATAATAAAGTGTGCACATCGCAATATTTTGTTTGGTACATGATCTTTCTACCATTTTACCTCTCAAGAACGCACATTGGTTGGAAGAAGGGGCTTTTAATGGCCACGCTTTGGGTAGGAACGCAGGGAATTTGGTTAAGCCAAGGTTACTATTTGGAATTCGAAGGCAAGAATGTAT tpg|BK006943.2|:459081-462067 7X173= 149=1X138=7X 
 tpg|BK006943.2| 177127 + tpg|BK006943.2| 177080 - INS TCAATAACGTGGATTTGAACTTTCAAAACACCTTTTATTTTCTCGATGATTTTGGACTTTTTTTTCTTTCCTAGCCTTGAGCCGTAAAGAGCGGAAAAACCATCAGACAATTCCAGAGCATTTTTTCTTTCTTGCGTTGTCAGCCCCGAACGTAAATAATTTCGAGGAGTCGATGGCCGTAGCAATAATCGAATAACACAATATATTGACGTCCACATCGCTTCACTTGCCGGTGCTTGAAATAACATCCCCTCAATACTCTGTCATAATT tpg|BK006943.2|:176524-177683 7X82=53S 5S1=174S 
 tpg|BK006943.2| 140304 + tpg|BK006943.2| 140386 - INS GGGCAATGCTGATGAGCAGTGAGCAGCTAGGATTCAATAAACGGGATTAACAAAAAATTGATATGTCCAAGCTTTCGAAAGATTACGTATCAGATTCAGACTCTGATGATGAAGTGATATCAAACGAGTTCAGCATACCAGATGGTTTCAAGAAATGTAAACATTTAAAGAATTTCCCTCTCAACGGTGATAACAAAAAAAAAGCGAAACAGCAACAGGTTTGGC tpg|BK006943.2|:139840-140850 7X6=19S 211=7X 
 tpg|BK006943.2| 131731 + tpg|BK006943.2| 131988 - INS TAAATATATTATAGAATCAGATCTGTGCATGAGTTGTTGCAAGAATTAAAGATATCATTGATACAACGAGAAACAAATTTAAACATTTGCTTTAAAAGATTGGAATAATGGGAAAGTAACGTCTTGTTATCGGGTCTTTTTTTCAAAAGGTACTCTTGTATCATACGGCATTTCCTCATCAGTTTCCAAAAATTTGTGATTATTGCTGGAAAAGTGTATTTAACATTGATGC tpg|BK006943.2|:131253-132466 7X6=226S 218=7X 
 tpg|BK006943.2| 43475 + tpg|BK006943.2| 42920 - INS GCACTACCTCAGCATTACGACGTGATGGATCTTTGCACTACCTCAGCCCACGCATCCAAAACGGCAAGTTCAATTTTTCTTTTCGCTTTGGGTGTAACGATTATAGCTTCCCCTATCCGTATACCGGAATTAGGATCTTTAAAGTTACCAAGAAGGTCAATTAGTAATTGTGAAATTCTTCCCAATTTATCTGGTGGCATTATATTCGATGCCAACACTTCAGCAGCAACAGTAATAGCAAAGGACATTACAGTAGGTGAGCTTCCTTTACTAAAAGCAGGCATTAATGCGCTAGTTATTTGGGCCTCTTGCTGTTCTAAAATCGACGATCCAGGAACCTGAGGATCTCTCATGGTGGAGTAGTTCTTGAGAACAAAATTCAAAATGTGTAGTCC tpg|BK006943.2|:42116-44279 7X7=312S 371=7X 
 tpg|BK006943.2| 402317 + tpg|BK006943.2| 402403 - INS TTTGGGTAAGACGCGAAAATGGAATATAATGACAATGTAAATATCGTCATCTTGAGATAATTATCAACAAGGTTGTCATGAGGAGTTACAGATAAAAGTCAACAGAGTGGAGTTAGTGGTGTTTTAACTGTAGTGCTCCATAGTTTCACGGCGGTTTCTCTTGTTTTCAGTTGGTAGTAACTTTTATCCTGGAAGTGCTGGAAATGAATAACTCAAATGAGCATAGGCG tpg|BK006943.2|:401845-402875 15S106= 68=54S 
 tpg|BK006943.2| 629628 + tpg|BK006943.2| 629406 - INS GTTTGAAAACAGCTTTTATGTCATATTCTTGAAATAGTTCACGCAATTTTCTCTTATCATTCTTTGGAAATTTAATCAAAGAAACCTTTGCGTTCTTTTCTTTGATGTGTTCCTGTAGATACGTTTTAGTGGTCTCATTAGTTGTGTATATTCTGTAACCAATAGTGGCCACTATGGAAGCCACTTGGCCCAAGTATTCTCGAGATGTATCACCTCCAAATAATATACCACTTGGAGGTAGTGGTACATGGAAGTTCATGGTAC tpg|BK006943.2|:628864-630170 7X243= 132=7X 
 tpg|BK006943.2| 554000 + tpg|BK006943.2| 554498 - INS TACGTGTAGCATTGATTTAGCTTCTGTTCATCATCATCTTCAGGATATCCTATTATAGTGTAGCATTGAAATTTCTCGGATATTGATTTAGCCAGTTCAAAAGAGGGCCCTTCATCTTTCTTAGTAACATAAGGTAAAATATCTTTTCTGGCATGAAAACTGTAACCTGTCAATGCAAATTCGGGGAATAGTATTACGTCTGGTTTCACATAGGTGGCACTTTTCGTAACTTTATCCAATATTGACCATGTTCTCTTAATTGTTTGATCTACTTGCCCAATTTGCGGATTGAGTTGAATTACTAGTACCTTTAGTGATACTAAAAGTTTTGTGCTCATCTTAGCACCATGAATTGCGTCTATTAGCATTCACTGAATGTCACGATAGAGTTATCGCTGTAAACTAGCACTTTTTAGCATTGAAATGCTTAAAATGTGTGAAACTAAAGTGGTTTTATTTCCAAAGAAGGGTTATCCCTTACTAGGGCAACGAATGAATATCTATTAGGGCTATAAAACAAAAATAGTTAAGTGAGATATATACCCTCTTGAATGGTGCAGGGT tpg|BK006943.2|:552860-555638 7X12=40S 179=1X366=7X 
 tpg|BK006943.2| 216739 + tpg|BK006943.2| 216144 - INS AATCAGTCTTCCTTATCTGAATGTTTTGCCTCTTTAGCATCTAAGTTTGAAAGAATGGTTTCCATGGCAGCTAAGATAATTGTTTTCTTTAAAGGCAAAGCTGTAGCAAATACAACTAATATGGTATGTGCAGCTATTTGACAATCCTTTGATTTAGAGGCTAAAAGTTTAGCAGATATTTCAAGTA tpg|BK006943.2|:215756-217127 7X178= 5S171=7X 
 tpg|BK006943.2| 637866 + tpg|BK006943.2| 637994 - INS ATCCAGTTCCACGCGATCCTATTTCTTTGCCTCTTGTTCAGAGGCACAGGAATGACAGAAGCCTTGGCCACGCCTGTGTTGAATGTCTTGGTCATCATCAGCGGAGCTAGTTCGTCGAGTGACTTTTCCAAAGCCTGGATGGGGTCCTGCCGGGTCTGGCAGTACACCAGATATAAGGC tpg|BK006943.2|:637494-638366 7X3=86S 85S5=7X 
 tpg|BK006943.2| 64973 + tpg|BK006943.2| 65660 - INS TGTCAGAGGGATCTGATATTGCCACAGATAGCAATGTTAGTACTTTTTTGAATTCTTCATATGAAATAACTCCGCTTCAATTTCTCGAACTACCGATAAAGAAACTACTAATACCAGACATGTTTGAAAACCGTTTAGACAAGATAACTTCAAATCCGAG tpg|BK006943.2|:64639-65994 191S12= 80=7X 
 tpg|BK006943.2| 127763 + tpg|BK006943.2| 127889 - INS CCAATCATGCCTAATTTATCCATACTTGGTAAGTTGCAATGGCTGCCAATACAAAAGACTGATAAGCATGGTAAAACGCCCGATTCTGATATCAAATCGTCATCCGTAATAAGGTTTAGTTTCTTCAGGAAGAAGTAAAATCTTCGTAACAGTATCGACC tpg|BK006943.2|:127429-128223 7X249= 80=7X 
 tpg|BK006943.2| 305382 + tpg|BK006943.2| 305526 - INS AACCATTTCATAGTTACACTTTAGGCGACTGATTTTTCATTAAATGGAAAATATCACAAGAAATTTCACGCTGGAGAAAAAAAAGGTTAGTCATCACTGATCTTCCCATGGAGTCATAAGCACGTTCGACATAAATTGTGAAAGTTAACACATTTGAAGCTAGGACCGTCAATCTAGGACACTAGTCGGTTACTTTTATCATGTGGAGGAGAATATTCGCGCATGAACTCAAGTATGATCAACCCAATGCATCTTCAAAAAACTTGATCC tpg|BK006943.2|:304828-306080 7X149=53S 3S1=220S 
 tpg|BK006943.2| 592552 + tpg|BK006943.2| 592557 - INS CTGTAAAGTTAGTCGCTCCAAATTCTTACATCCGACAAAATAGTTAAGCTCTGTATCGTGCATGTAGTCACCAACAAATGAAAAATTTAATCTTTTGATCATTAAACGATAGTTGAATACAGTTTCTTCAGAAGTTAACTTCATAGTCCTTAAAAACAAGTCTAATTGACTCTTTTTGTTGATGTGCGGTCTGTAATAAAG tpg|BK006943.2|:592136-592973 7X6=94S 95S6=7X 
 tpg|BK006943.2| 589212 + tpg|BK006943.2| 589300 - INS CTCCAGATAGGCAATAGCAAAACAGCCAGCATTCCCGCTGATATTCATCCTAAACCAAGGAAAAACTTGCAAGAACCAAGAAGCCTATCAATAAGTGGAAAAGTTGTTCCAACAGAAAGAAAATTAGATAACATCAATATAGATCTAAATTTTTCGGCGTCCGATTTTTCACCATCATCACAATCTGAGCAATCATCAAAAAGCTCAAGCGTTATTTCAACGCCGGTAGCGAGCCCTAAAATTAATCTCACACGCAGTTTGCATGCAGTCAAAG tpg|BK006943.2|:588650-589862 7X253= 7=1X249=7X 
 tpg|BK006943.2| 27360 + tpg|BK006943.2| 27437 - INS GGGAAGCTTGGCGTGTTCCGCTTGGTCTATGTTTTGCATGGGCTATTATTATGATTGGTGGTATGACGTTTGTTCCGGAATCTCCTCGGTTTTTGGTGCAAGTCGGTAAGATTGAGCAAGCTAAAGCTTCTTTTGCCAAGTCGAACAAGCTTAGTGTTGACGATCCTGCTGTGGTTGCAGAGATTGATC tpg|BK006943.2|:26968-27829 7X4=159S 178=7X 
 tpg|BK006943.2| 365866 + tpg|BK006943.2| 366160 - INS CCCTACCACTGATCCGATATCCACAGGCTCCAATACTTCTAGAACGAACGATAATGCTCATATTCCTCCGACCGATGCGCCTGGATTTGATAAATTTATGAACAATGCAGAGGAAAATGCCATTGACGCTGCTTATGATGATGTGCTAGACAAAATCCAGGATGCG tpg|BK006943.2|:365520-366506 7X4=79S 78S5=7X 
 tpg|BK006943.2| 129180 + tpg|BK006943.2| 129169 - INS ATTACATTATCACGTACATAAAAAACCATCAATGCTACGTTTCCTGATCTTTTCGTACATAAAAGATTGTGCGTATCAGCCACAAGTAAGCTTGGACTTAAGATACACAAAAATAAAAAGTAAAATTTAAAATTTGTCTTCCAAAGGAGAGTCATTGAGCAGTTGATGAAGTTTAGTTGAGCTTTGAGAAAGCTCACCTACTTGGCTTGTACCCTTCTCTTTATATGTACTCACTGCAGGGATGTTTGCTTTAATTTTGGTGACCTTTGTGCCATAGGCCCTAGGCTCCAGCTTGATCAATGTGTGTAGTGGGATTGACATCCAAGG tpg|BK006943.2|:128501-129848 7X110=1D99=2S 307=7X 
 tpg|BK006943.2| 390902 + tpg|BK006943.2| 391045 - INS AACCTCCTTAATTTCTTTATCTTTTTTTCCCTTCACCTCTGTGCTCTTTTTTTAGCCACAGCTGTGCATTACGCTTGCTTTGCTTGTTTTGTTCTCTTTCGCCATGCCATATTACTACTTTTCTACTTACTGGCACGAGGCCGCGCAAGCCAGATCCAAGCACGCCAGAAAGTGCGGTGTACTGGTG tpg|BK006943.2|:390514-391433 7X42=51S 2S1=166S 
 tpg|BK006943.2| 607294 + tpg|BK006943.2| 607456 - INS ATGCAGGACGGGCCGTGGCGGAAAGAACAGCATGATATAGATAATATATGATATGAATTGATTTTTTTTTCTTTTTTTCTTGCGGCTGGTATGGTATTGTAAGGATGATAGTGCATTCTATGAGTGATTTTTGTGACGGTGACGTACGATCTCTATACCTT tpg|BK006943.2|:606958-607792 7X9=71S 77S4=7X 
 tpg|BK006943.2| 377151 + tpg|BK006943.2| 377639 - INS CGTCAGTTTCTCAAGCTGACACTTGATTTATTCTAAACAAATTTCAATCTTGGACAATTAGTTGACATAAACTACGTTACTAATTTTTGTTGTATTAAGGGCTTAAATAATACCGGATGTCTTGGCAATTCTATCGTTAGGAGAGTAATAGTTGTCAGACTTATTGTCGGCTTGTTCGCACATCGTTACTTATCCTATATTATAC tpg|BK006943.2|:376727-378063 7X137=16S 3S1=161S 
 tpg|BK006943.2| 723956 + tpg|BK006943.2| 723237 - INS CCACATCTTAATTCAAGGATGTACTGTTTATAATCAGGATGACTGTATTGCTGTGAATTCCGGTTCAACTATTAAATTTATGAACAACTACTGCTACAATGGCCATGGTATTTCTGTAGGTTCTGTTGGTGGCCGTTCTGATAATACAGTCAATGGTTTCTGGGCTGAAAATAACCATGTTATCAACTCTGACAACGGGTTGAGA tpg|BK006943.2|:722813-724380 7X6=242S 103=7X 
 tpg|BK006943.2| 719798 + tpg|BK006943.2| 719607 - INS CTGACTTCAATGTTGTTATGTTAAACACATTGAAGAAAACAACAAAACAAGGATAATCAAATAGTGTAAAAAAAAAAATTCAAGATGTCAGCGGATGCTAGTACAAATTCGAATGCTTCCCTAGACGAAAAAAATTTAAACATCACTTCAGAAGCTGAAATCAAGAATGAAGACGTAACCGCGGAGCCAGTTCTAAGCACGGTACTATCACCCAACGGTAAAATTGTCTACATCAGTGACAAGGTTGATGAGGCCATGAAGTTGGCTGAAGAAGCCAAAGAAATCGAAGTGACACCAGAAGAAGATAGAAAACTTCGTTGGAAGATCGACTATTGTATGTTTCCTTTGATGTGTATATTGTATGCTGTTCAATTTATGGACAAGATTTCCACTAGTTCAGCGGCGGTCATGGGATTAAGAAC tpg|BK006943.2|:718749-720656 7X237= 13S396=7X 
 tpg|BK006943.2| 553135 + tpg|BK006943.2| 553334 - INS TTAAATTCTTGCCTTCGGAATAGGATAATAACAAAAACCATTATTTATTCATTCTTGCCTCACTTAAATTCGGCCCTTACGGCGACATTTCAATAACATAAATATGCGTGTAACCTTATTAATTTATAATGTCTAATTTATTATAATATTCCTTCACCTAAACACTTCAAATTGGACCTCACGCAATATAGCGC tpg|BK006943.2|:552733-553736 7X255= 182=7X 
 tpg|BK006943.2| 104364 + tpg|BK006943.2| 105045 - INS CTTTTGAAATCTCACTTCAGAAACGAAAAATACTACATAGATATCACCGAATTGTTCCATGAGGTCACCTTCCAAACCGAATTGGGCCAATTGATGGACTTAATCACTGCACCTGAAGACAAAGTCGACTTGAGTAAGTTCTCCCTAAAGAAGCACTCCTTCATAGTTACTTTCAAGAC tpg|BK006943.2|:103992-105417 7X13=76S 84S6=7X 
 tpg|BK006943.2| 313566 + tpg|BK006943.2| 312856 - INS GGGAGACCAGAGTGAACGAAAGTGCTGACAAAGTAATAGGAGTGATCAAAGCCGTGAACTTTTTTTATTTCCACGTAGTCCTGCCATGAAGTGGCTTTCACCGCCTCAAGTAGTAATTCCGGTTTCAAGTGTTCTTCCAAAAAGGGATCGGAGTCTCCTACAT tpg|BK006943.2|:312516-313906 7X5=5S 3S150=7X 
 tpg|BK006943.2| 217397 + tpg|BK006943.2| 217747 - INS GTCAAAGTTACACAAAGAGTGAAGAAGCAAATAGTCCCACAGAAATACCGACACAAACTTGAATCATTGTCATACCAAATGACATTGAGGACGATGGATCGGAGGTGCTTGTCGTAATGGTTTCATTAGCATTAACAATTGTATTTGCACTTTGCAACCCAGACAACAACGAATTTTGTGAAGCAATACCAGATGGCACTTGAACGAAGATTGCGGGAAGCATAGCTGATACCGCTAAACCTTTCCAAATTCTGGAATATAGATTACCTAAAAC tpg|BK006943.2|:216835-218309 7X161= 257=7X 
 tpg|BK006943.2| 259786 + tpg|BK006943.2| 260185 - INS GGTCTTGAGTGGCCGGTAGTTTTTATTCCTGGATGCGAAGAAGGTATAATTCCTTGTGTGTTCAACGATGATAAGAAAGACGAATCAGAGGAGGACGAAGAAGAAGATCAAGAAAATAGTAAGAAAGATGCAAGCCCAAAAAAGACTAGAGTTTTATCCGTGGAAGATTCTATAGATGAGGAAAGAAGAATGTT tpg|BK006943.2|:259384-260587 7X5=337S 97=7X 
 tpg|BK006943.2| 617003 + tpg|BK006943.2| 617149 - INS CAAACTTGAATGAAGTATATAACGAAGTCAATGAAACCTCTCCCATACTAGGTTCGGAACCTGTTAAGGGGAACAAGACCGCGCACTTGTTATGAAAATTCTTCCTATAACTATATTGAAAGCTATTTTTCCACATCGGCAGACAAACGACTGTCC tpg|BK006943.2|:616677-617475 7X48=30S 1S1=23S 
 tpg|BK006943.2| 380990 + tpg|BK006943.2| 381666 - INS TTAATATGCTGCTACTCTCCGTGGTCGACATTAAGAGATTGATCGGTTTGAAATATAACGACAGATCTGTTCAGA tpg|BK006943.2|:380826-381830 7X7=12S 6S51=7X 
 tpg|BK006943.2| 428688 + tpg|BK006943.2| 428657 - INS GTACCTCTCCGGTGATACAGTTTTGAAATGGAGCTCTTTAAAGACTTTAATGTTGAATAGTAACCAAATGTTATCTCTGCCTGCAGAATTATCAAATCTCTCACAGCTAAGTGTATTTGATGTTGGAGCAAATCAATTAAAGTATAATATATCAAACTATCATTACGATTGGAACTGGAGGAATAATAAAGAACTAAAATATTTGAATTTTTCAGGAAATCGAAGGTTTGAAATAAAGTCATTTATAAGTCACGATATTGATGCTGATTTGTCAGATCTGACAGTATTACCTCAGTTAAAGG tpg|BK006943.2|:428039-429306 7X269= 284=7X 
 tpg|BK006943.2| 80507 + tpg|BK006943.2| 80540 - INS CAACTAAAGGATCAACACGGCTTTAAAGTGTTTTATATATACGCAGATATGAAAAAAGCATTTTCACGGTTATTGGAAATTTTTATTTTACGACTGGTTCCTAGCACAACAAGAGGATATACTAATAGTTCAGGTTACAATGCTGATTAGGTTAAAGAAGAGAA tpg|BK006943.2|:80165-80882 7X4=78S 68S14=7X 
 tpg|BK006943.2| 646026 + tpg|BK006943.2| 646291 - INS CCTTTTAATATGATCTAGAGGTAAAATTGACTAAGTAGTCAGATCTTATTCTACATTGAGCCTGCGTTGTCAACATGCACATCTCTGTCTCTTGGGATGATAATTTTTCAATGATGATTCCAGGGTTACTTTAACGTTACACAAAAGAAATTAATTAGTGCGGCTGTTTCTGTGAGCGGGGCAGTAAGTCCGAAGCCCTTGATATTAGCCCATACCCTACACATTTTACTCGTTTGCCCTACATCAGATAAAATACTGGCCCTAAGCCCTCCTAATCTCTTCTGGTT tpg|BK006943.2|:645438-646879 7X100= 144=7X 
 tpg|BK006943.2| 100382 + tpg|BK006943.2| 100717 - INS CTTTACCCACTTCGCAAGTACACGATTCATTGTTGGTGATATCTTTAAACTTATTCACATCTACGTAGGAGCCTGTAAAACCAACATTAGTGAAATCCAACTTTTGGTACGACTGAGGTCCACTGGCAGCGACTGTGTGCAACATAAACATGCACACGGAAAGGACTATACTCTGTAACATTTGTCTTATTTAAGCTTGTAATGTTTGCACTTGAGTATGTTCTAT tpg|BK006943.2|:99916-101183 7X172=1X57= 113=7X 
 tpg|BK006943.2| 300154 + tpg|BK006943.2| 300557 - INS TGTAGTTTAGCGA tpg|BK006943.2|:300114-300597 7X6= 4S3=7X 
 tpg|BK006943.2| 68868 + tpg|BK006943.2| 69023 - INS TGCGCTGCACTATTTTCATCAATAGTACCATATACGTTCATGTCAGCTATACCAATAACTCCAACTAAGCGTATCAGAAGAAATCTATTTGACGATGCTCCAGCAACGCCTCCACGACCTTTGAAAAGAAAAAAGTTGCAGTTCACAGATGTTACACCAGAATCATCC tpg|BK006943.2|:68518-69373 7X75=51S 7S1=149S 
 tpg|BK006943.2| 437612 + tpg|BK006943.2| 437142 - INS GTTATTCTGTATCAGTAACTTTAAATAATGCTGGTCGCCCGCGCATTACTAATTTGGCTAACAACGATAGAGTTAGTACAGCCAGCATGGCTATTCACGATGATGATTATGGGTCCATCCAAAATTCAACAATTGGGGATTCTGGGTCAATATTACGCCCTACTGCCTCCTTAACAGAAATGATGAGTGGTGGAGCGGGGAGAAGGTTTACAAATAATGACATGGATTCAATTGTAG tpg|BK006943.2|:436654-438100 7X4=230S 223=7X 
 tpg|BK006943.2| 191377 + tpg|BK006943.2| 191416 - INS GCCTTGGATTCTTTCTATTAGAAAAGCAGAGAATAAATAGACATGATACCTCGCCTTCTATCCTCTGCAGCGTATTATTGTTTATTCCACGCAGGCATCGGTCGTTGGCTGTTGTTATGTCTCAGATAAGCGCGTTTGTTATGCGAAAAAAAAAAACTTTACAGAGGCTTTGTTTATATATAGAAAGACCACGAAAAAAACAGTGATGGCTTCATGCTTTTCAGTTTCATTATTGGCACGAGTAGCAGTCGTTGAGCCCATCAGAGTGC tpg|BK006943.2|:190825-191968 7X7=29S 36=1X1=1X2=1X211=7X 
 tpg|BK006943.2| 458373 + tpg|BK006943.2| 459108 - INS ATCCTTAGAGCTATCCTTAAATCGTAAACTAGTTCACAAATATCACTCTTTAGTGCAAGG tpg|BK006943.2|:458239-459242 7X11=26S 13=1X31=7X 
 tpg|BK006943.2| 268112 + tpg|BK006943.2| 268301 - INS GCTCTTCCTAGAAATTCCTTT tpg|BK006943.2|:268056-268357 7X3=7S 11=7X 
 tpg|BK006943.2| 92933 + tpg|BK006943.2| 93120 - INS CAGTGGTACTGGTTTTCTTTGGATTGGCACTTTTGGAGTGATCGTTCATGATTTCACGTTCCTGTTCGTTTCTCTCTTCGCCACTATCTACCTTCTTATCTACACTTTCCGTCTTTTCTATGATATCCTCCTGTTCAGCTTTATGCGCATCTGGAATTTCAGATGGAGTATTAGCAACCGACGAAGTGTTGCCT tpg|BK006943.2|:92531-93522 7X12=85S 92S5=7X 
 tpg|BK006943.2| 397965 + tpg|BK006943.2| 397995 - INS ACCAATGAGATCTGTTAAGAAGTATTGTGGAGAATATCTTCATGATTTGGTTTTTCTATTAACCTTCTTAATCTTTTCTTTCTTCATCTGCCATCGCCTTTCTATGTTTTCCGTATTTCTTCCCCGCAAGTTCTTTAAACTCAGATAGTATTAGAATCGATAATTAAGGCCAGGTCAAAGTTCGTATTAATTTCAACCTTTGGGCACCTATAT tpg|BK006943.2|:397525-398435 32S55=26S 103S4=7X 
 tpg|BK006943.2| 683553 + tpg|BK006943.2| 683805 - INS TTTTTCCGAAAATATGGCTAGCCAACTTAGGTGAATGGGGAAGGGTACTAGATTCATTCATTTATTTCTATTCAAGGACAAGAACTTTTAACATAGTAAGACCTTTATGTTAGTTTGGTGCGGCTGACAAATTCATAGCTAATGTGCTAGAGCTCTTATAT tpg|BK006943.2|:683217-684141 7X6=74S 75S6=7X 
 tpg|BK006943.2| 262070 + tpg|BK006943.2| 261866 - INS ATCCTACAAGGTAACAGTATTAGCGTGTTTAGAAGGTATGGTTCACTAGCATAAATAGTAATAGATAGAAGCAAAGCAACCCAGTTCAATGCAAAATCAATTATGTATTGCACGCTGGAAATGCCAGGAGGCATAAGGTTGGAATTTTTCAATAAGTTCCATGA tpg|BK006943.2|:261524-262412 12S124=15S 15S5=7X 
 tpg|BK006943.2| 56319 + tpg|BK006943.2| 56308 - INS CGACAACAAAATAGCTTATGACTATTAAATCGGACTCTTAATTTTTAGCTAATATCTCTTCAGAATTTATTCGTTTCTTCGTATATTACCAATATAATTGATTGCTGAACCAGCTTTGAAAAAATCGATTTGATCTTTAGACATAGTATGTTTTGCCTTGATGGTGAACGATTCACCGTTTGGTTTAGTAATTTTAACATCAATTTCACCACCGTTATTACCATCCTTAGCAATCATGTCAACTAGGTTCAACGTTTCTAAAACATCTCCGC tpg|BK006943.2|:55750-56877 7X14= 255=7X 
 tpg|BK006943.2| 328554 + tpg|BK006943.2| 329146 - INS ATCCATTTCTGGAATAAAGTATTTGTTTTTGCTGAACTGTCCCTGCTTATTGTTACTATCGTTTTGTAGGGCGTAGTGCCGATGATTTCTTTCCAATGACTGAAAATATCTTCTTGAAAAGCTTGAATTGGCAAATTCAAATCCAAGTGGCACAGTGTTCTCTGGAATACTGAGCCTACTGCTTTCTGATTCTACTCCAGCAGAGGCTCGACGATGAAGTTGTCTTCTGTTTATAATATCAGGGTTAATTTCCGTACCACAT tpg|BK006943.2|:328016-329684 14S45=79S 125S6=7X 
 tpg|BK006943.2| 386848 + tpg|BK006943.2| 386641 - INS TTCTGATGTTTTCTTCAGAGCTTCAATTGAGTAAATTTTTTCATCTCTCATATTCAAAACATTTTCAGTCAAGCTTCTATAATCATATATTTTCTTTTCGTCTTGAACTCTCTTTTGTCTCAGTAATTCCTTGGTCCACTGTTTCCTTTTAATGCCATGCTGTTTAATG tpg|BK006943.2|:386289-387200 7X11=73S 78S7=7X 
 tpg|BK006943.2| 580705 + tpg|BK006943.2| 581015 - INS AAACAATGAAGATTTGAATGAACGAAATTTAATCAGGTTTGACCAAAAATTCAGCCATTTATAGGAAAGGGATAAATGGTTCAAATTGTGAATGGAAACTAGGCAATCCTTTTTGATACAAATTGGAATATCTGGTTGAACAGTGATAGATGCAATTTTACCATTTTCGTCTACTAGCCTGAAACGGGAAGTCGCAATATCCTTGCTTAAGTTCTCGATATATGTCCTTTCTTTAGTTACGACATTAC tpg|BK006943.2|:580195-581525 7X232= 16S5X2S 
 tpg|BK006943.2| 645276 + tpg|BK006943.2| 644895 - INS AAGTATTTAACGTGATAATATAGTC tpg|BK006943.2|:644831-645340 7X4=8S 10=1X2=7X 
 tpg|BK006943.2| 167763 + tpg|BK006943.2| 167945 - INS GGAGGTTAGTAACCAACGGAACCGAATAATCGACAGCCAAACGACG tpg|BK006943.2|:167657-168051 7X3=14S 23=7X 
 tpg|BK006943.2| 89017 + tpg|BK006943.2| 89320 - INS CAATAGCCTAAGATTCTCGAAACCACTTCCTTGCAGAATTCAGGTAAGGAAGTGAGAAATTGAGTAGAACGTTGAATGAACTCAGCACGGAAATCTTGAAAAGAGCCTCCTCTGGTATTCAAGAATGATACAACCATCAGGTATATCAATGTAAACAGTAGAGCGTATAGGAATAACCAAGTGAACCACGAAGTCCCGCCTGCCTTCTTAGCTGGCTTTTTCCCCTCGCTGTCAC tpg|BK006943.2|:88533-89804 12S112= 118=7X 
 ref|NC_001224| 78660 + ref|NC_001224| 79190 - INS GGATAATATATATTATTATAAGATATATATATAACAATAAATTTATGACACATTTAGAAAGAAGTAGACATCAACAACATCCATTTCATATGGTTATGCCTTCACCATGACCTATTGTAGTATCATTTGCATTATTATCATTAGCATTATCACTAGCATTAACAATGCATGGTTATATTGGTAATATGAATATGGTATATTTAGCATTATTTGTATTATTAACAAGTTCTATTTTATGATTTAGAGATATTGTAGCTGAAGCTACATATTTAGGTGATCATACTATAGCAGTAAGAAAAGGTATTAATTTAGGTTTCTTAATGTTTGTATTATCTGAAGTATTAATCTTTGCTGGTTTATTCTGAGCTTATTTCCATTCAGCTATGAGTCCTGATGTACTATTAGGTGCATGTTGACCACCCGTAGGTATTGAAGCTGTACAACCT ref|NC_001224|:77754-80096 22S7=1X9=223S 9S424=7X 
 ref|NC_001224| 11141 + ref|NC_001224| 10891 - INS AGATAAATATATTTATAGTGAATACCTTTTTTAATATTTATTTTTAATATTTATTTTTAATATTTTATTTTTAATAAAATATAATCTTGTAAGTAAGAAAAGAATTTCGGTGATTGGAACCTTGAAAGGATAAATTTCTTATTTATTATAATATTTATATTAATAGTTCCGGGGCCCGGCCACGGGAGCCGGAACCCCGAAAGGAGTATTATTAAACATTTAATATATTATATTAATATTTAATTTAAATG ref|NC_001224|:10375-11657 13S112=1X6=53S 126=7X 
 ref|NC_001224| 52189 + ref|NC_001224| 52190 - INS CCCTATTATTATATATAATATAAATATTTATATATTATTTTTATATTAATATTTATAGATGGGGGGTCCCTATTATTATTGAAAATAATAATTATTAATGGACCCCAGATAGCTTCTTGTTTATCATTTATATATATATATATATTATTAATTATTTTATTCTCCTTTCGGGGTTCCGGCTCCCGTGGCCGGGCCCCGGAACTTTATAATATTATTATTAATTATTTAATTAATATTATAATCATATAATTTAATATTTTATTTAATTTTATTAAAATTTAATAT ref|NC_001224|:51605-52774 7X23= 3S265=7X 
