 tpg|BK006942.2| 44338 + tpg|BK006942.2| 44631 - INS 
 tpg|BK006942.2| 122627 + tpg|BK006942.2| 123122 - INS 
 tpg|BK006942.2| 388041 + tpg|BK006942.2| 387330 - INS 
 tpg|BK006942.2| 249460 + tpg|BK006942.2| 249837 - INS 
 tpg|BK006942.2| 86083 + tpg|BK006942.2| 85775 - INS 
 tpg|BK006942.2| 390815 + tpg|BK006942.2| 390625 - INS 
 tpg|BK006942.2| 311882 + tpg|BK006942.2| 311131 - INS 
 tpg|BK006942.2| 151450 + tpg|BK006942.2| 150734 - INS 
 tpg|BK006942.2| 408273 + tpg|BK006942.2| 408538 - INS 
 tpg|BK006942.2| 283628 + tpg|BK006942.2| 284122 - INS 
 tpg|BK006942.2| 380541 + tpg|BK006942.2| 380383 - INS 
 tpg|BK006942.2| 215400 + tpg|BK006942.2| 214804 - INS 
 tpg|BK006942.2| 330980 + tpg|BK006942.2| 330206 - INS 
 tpg|BK006942.2| 404602 + tpg|BK006942.2| 404560 - INS 
 tpg|BK006942.2| 105552 + tpg|BK006942.2| 105876 - INS 
 tpg|BK006942.2| 94080 + tpg|BK006942.2| 93935 - INS 
 tpg|BK006942.2| 50128 + tpg|BK006942.2| 50576 - INS 
 tpg|BK006942.2| 247102 + tpg|BK006942.2| 246544 - INS 
 tpg|BK006942.2| 334228 + tpg|BK006942.2| 334000 - INS 
 tpg|BK006942.2| 254258 + tpg|BK006942.2| 254193 - INS 
 tpg|BK006942.2| 415987 + tpg|BK006942.2| 415739 - INS 
 tpg|BK006942.2| 196605 + tpg|BK006942.2| 197062 - INS 
 tpg|BK006942.2| 269061 + tpg|BK006942.2| 268770 - INS 
 tpg|BK006942.2| 56274 + tpg|BK006942.2| 55664 - INS 
 tpg|BK006942.2| 48662 + tpg|BK006942.2| 49293 - INS 
 tpg|BK006942.2| 200673 + tpg|BK006942.2| 199993 - INS 
 tpg|BK006942.2| 384860 + tpg|BK006942.2| 384686 - INS 
 tpg|BK006942.2| 84780 + tpg|BK006942.2| 84304 - INS 
 tpg|BK006942.2| 73802 + tpg|BK006942.2| 73195 - INS 
 tpg|BK006942.2| 279127 + tpg|BK006942.2| 279648 - INS 
 tpg|BK006942.2| 92636 + tpg|BK006942.2| 92434 - INS 
 tpg|BK006942.2| 434688 + tpg|BK006942.2| 434441 - INS 
 tpg|BK006942.2| 403464 + tpg|BK006942.2| 403040 - INS 
 tpg|BK006942.2| 414244 + tpg|BK006942.2| 413660 - INS 
 tpg|BK006942.2| 222005 + tpg|BK006942.2| 221726 - INS 
 tpg|BK006942.2| 243836 + tpg|BK006942.2| 244571 - INS 
 tpg|BK006942.2| 36723 + tpg|BK006942.2| 36440 - INS 
 tpg|BK006942.2| 322441 + tpg|BK006942.2| 322269 - INS 
 tpg|BK006942.2| 127355 + tpg|BK006942.2| 126800 - INS 
 tpg|BK006942.2| 67272 + tpg|BK006942.2| 67163 - INS 
 tpg|BK006942.2| 162865 + tpg|BK006942.2| 162388 - INS 
 tpg|BK006942.2| 280850 + tpg|BK006942.2| 281081 - INS 
 tpg|BK006942.2| 216661 + tpg|BK006942.2| 216844 - INS 
 tpg|BK006942.2| 57249 + tpg|BK006942.2| 56483 - INS 
 tpg|BK006942.2| 397299 + tpg|BK006942.2| 397118 - INS 
 tpg|BK006942.2| 220895 + tpg|BK006942.2| 221141 - INS 
 tpg|BK006942.2| 37316 + tpg|BK006942.2| 37199 - INS 
 tpg|BK006942.2| 342744 + tpg|BK006942.2| 342885 - INS 
 tpg|BK006942.2| 153082 + tpg|BK006942.2| 152537 - INS 
 tpg|BK006942.2| 400770 + tpg|BK006942.2| 400764 - INS 
 tpg|BK006942.2| 368855 + tpg|BK006942.2| 368933 - INS 
 tpg|BK006942.2| 183657 + tpg|BK006942.2| 183641 - INS GCTA
 tpg|BK006942.2| 356842 + tpg|BK006942.2| 356243 - INS 
 tpg|BK006942.2| 103417 + tpg|BK006942.2| 103163 - INS 
 tpg|BK006942.2| 89059 + tpg|BK006942.2| 88460 - INS 
 tpg|BK006942.2| 163901 + tpg|BK006942.2| 164288 - INS 
 tpg|BK006942.2| 303613 + tpg|BK006942.2| 303122 - INS 
 tpg|BK006942.2| 52505 + tpg|BK006942.2| 52446 - INS 
 tpg|BK006942.2| 111902 + tpg|BK006942.2| 111381 - INS 
 tpg|BK006942.2| 335479 + tpg|BK006942.2| 334707 - INS 
 tpg|BK006942.2| 51522 + tpg|BK006942.2| 51715 - INS 
 tpg|BK006942.2| 353945 + tpg|BK006942.2| 353679 - INS 
 tpg|BK006942.2| 41391 + tpg|BK006942.2| 40823 - INS 
 tpg|BK006942.2| 231415 + tpg|BK006942.2| 231178 - INS 
 tpg|BK006942.2| 424002 + tpg|BK006942.2| 424744 - INS 
 tpg|BK006942.2| 290175 + tpg|BK006942.2| 290565 - INS 
 tpg|BK006942.2| 266454 + tpg|BK006942.2| 266449 - INS 
 tpg|BK006942.2| 361139 + tpg|BK006942.2| 360815 - INS 
 tpg|BK006942.2| 116903 + tpg|BK006942.2| 117644 - INS 
 tpg|BK006942.2| 187465 + tpg|BK006942.2| 187801 - INS 
 tpg|BK006942.2| 276441 + tpg|BK006942.2| 276622 - INS 
 tpg|BK006942.2| 382335 + tpg|BK006942.2| 382573 - INS 
 tpg|BK006942.2| 271521 + tpg|BK006942.2| 272141 - INS 
 tpg|BK006942.2| 82573 + tpg|BK006942.2| 82096 - INS 
 tpg|BK006942.2| 143638 + tpg|BK006942.2| 143275 - INS TTCTTCCACCA
 tpg|BK006942.2| 210830 + tpg|BK006942.2| 210945 - INS 
 tpg|BK006942.2| 212663 + tpg|BK006942.2| 212678 - INS 
 tpg|BK006942.2| 267460 + tpg|BK006942.2| 267584 - INS 
 tpg|BK006942.2| 323110 + tpg|BK006942.2| 323298 - INS 
 tpg|BK006942.2| 410490 + tpg|BK006942.2| 409786 - INS 
 tpg|BK006942.2| 115399 + tpg|BK006942.2| 116083 - INS 
 tpg|BK006942.2| 114014 + tpg|BK006942.2| 113941 - INS 
 tpg|BK006942.2| 393176 + tpg|BK006942.2| 393205 - INS 
 tpg|BK006942.2| 85182 + tpg|BK006942.2| 85025 - INS 
 tpg|BK006942.2| 224318 + tpg|BK006942.2| 224453 - INS 
 tpg|BK006942.2| 419964 + tpg|BK006942.2| 419339 - INS 
 tpg|BK006942.2| 233307 + tpg|BK006942.2| 233160 - INS 
 tpg|BK006942.2| 389174 + tpg|BK006942.2| 389879 - INS 
 tpg|BK006942.2| 121814 + tpg|BK006942.2| 121199 - INS 
 tpg|BK006942.2| 437262 + tpg|BK006942.2| 437514 - INS 
 tpg|BK006942.2| 195725 + tpg|BK006942.2| 196067 - INS 
 tpg|BK006942.2| 226472 + tpg|BK006942.2| 225843 - INS 
 tpg|BK006942.2| 126566 + tpg|BK006942.2| 126207 - INS 
 tpg|BK006942.2| 337695 + tpg|BK006942.2| 337157 - INS 
 tpg|BK006942.2| 341970 + tpg|BK006942.2| 341376 - INS 
 tpg|BK006942.2| 166219 + tpg|BK006942.2| 166109 - INS 
 tpg|BK006942.2| 136369 + tpg|BK006942.2| 136727 - INS 
 tpg|BK006942.2| 227469 + tpg|BK006942.2| 227852 - INS 
 tpg|BK006942.2| 80739 + tpg|BK006942.2| 80415 - INS 
 tpg|BK006942.2| 70195 + tpg|BK006942.2| 70141 - INS 
 tpg|BK006942.2| 148017 + tpg|BK006942.2| 148723 - INS 
 tpg|BK006942.2| 167204 + tpg|BK006942.2| 167767 - INS 
 tpg|BK006942.2| 422685 + tpg|BK006942.2| 423444 - INS 
 tpg|BK006942.2| 155345 + tpg|BK006942.2| 156007 - INS 
 tpg|BK006942.2| 169452 + tpg|BK006942.2| 169310 - INS 
 tpg|BK006942.2| 366884 + tpg|BK006942.2| 366727 - INS 
 tpg|BK006942.2| 176366 + tpg|BK006942.2| 175865 - INS 
 tpg|BK006942.2| 43801 + tpg|BK006942.2| 43844 - INS 
 tpg|BK006942.2| 256722 + tpg|BK006942.2| 257110 - INS 
 tpg|BK006942.2| 383877 + tpg|BK006942.2| 383117 - INS 
 tpg|BK006942.2| 91314 + tpg|BK006942.2| 90585 - INS 
 tpg|BK006942.2| 79647 + tpg|BK006942.2| 79163 - INS 
 tpg|BK006942.2| 394355 + tpg|BK006942.2| 394889 - INS 
 tpg|BK006942.2| 327249 + tpg|BK006942.2| 326852 - INS 
 tpg|BK006942.2| 309934 + tpg|BK006942.2| 309237 - INS 
 tpg|BK006942.2| 379396 + tpg|BK006942.2| 378636 - INS 
 tpg|BK006942.2| 61035 + tpg|BK006942.2| 60408 - INS 
 tpg|BK006942.2| 351640 + tpg|BK006942.2| 352061 - INS 
 tpg|BK006942.2| 373703 + tpg|BK006942.2| 373362 - INS 
 tpg|BK006942.2| 320968 + tpg|BK006942.2| 320367 - INS 
 tpg|BK006942.2| 273597 + tpg|BK006942.2| 273472 - INS 
 tpg|BK006942.2| 154647 + tpg|BK006942.2| 155056 - INS 
 tpg|BK006942.2| 247775 + tpg|BK006942.2| 247107 - INS 
 tpg|BK006942.2| 20067 + tpg|BK006942.2| 19452 - INS 
 tpg|BK006942.2| 77481 + tpg|BK006942.2| 78057 - INS 
 tpg|BK006942.2| 328795 + tpg|BK006942.2| 328123 - INS 
 tpg|BK006942.2| 299383 + tpg|BK006942.2| 298893 - INS 
 tpg|BK006942.2| 365105 + tpg|BK006942.2| 365832 - INS 
 tpg|BK006942.2| 125202 + tpg|BK006942.2| 125626 - INS 
 tpg|BK006942.2| 270722 + tpg|BK006942.2| 271020 - INS 
 tpg|BK006942.2| 364534 + tpg|BK006942.2| 365226 - INS 
 tpg|BK006942.2| 285787 + tpg|BK006942.2| 285076 - INS 
 tpg|BK006942.2| 71006 + tpg|BK006942.2| 71272 - INS 
 tpg|BK006942.2| 343900 + tpg|BK006942.2| 343986 - INS 
 tpg|BK006942.2| 406270 + tpg|BK006942.2| 405600 - INS 
 tpg|BK006942.2| 54186 + tpg|BK006942.2| 53892 - INS 
 tpg|BK006942.2| 53691 + tpg|BK006942.2| 53399 - INS 
 tpg|BK006942.2| 47634 + tpg|BK006942.2| 46955 - INS 
 tpg|BK006942.2| 282103 + tpg|BK006942.2| 282719 - INS 
 tpg|BK006942.2| 28823 + tpg|BK006942.2| 28932 - INS 
 tpg|BK006942.2| 127953 + tpg|BK006942.2| 128563 - INS 
 tpg|BK006942.2| 376094 + tpg|BK006942.2| 376558 - INS 
 tpg|BK006942.2| 300015 + tpg|BK006942.2| 299581 - INS 
 tpg|BK006942.2| 314889 + tpg|BK006942.2| 315556 - INS 
 tpg|BK006942.2| 259710 + tpg|BK006942.2| 259256 - INS 
 tpg|BK006942.2| 165538 + tpg|BK006942.2| 165250 - INS 
 tpg|BK006942.2| 162014 + tpg|BK006942.2| 161595 - INS 
 tpg|BK006942.2| 357602 + tpg|BK006942.2| 358062 - INS 
 tpg|BK006942.2| 201078 + tpg|BK006942.2| 201731 - INS 
 tpg|BK006942.2| 160653 + tpg|BK006942.2| 160843 - INS 
 tpg|BK006942.2| 245651 + tpg|BK006942.2| 245394 - INS 
 tpg|BK006942.2| 350231 + tpg|BK006942.2| 349890 - INS 
 tpg|BK006942.2| 212191 + tpg|BK006942.2| 211809 - INS 
 tpg|BK006942.2| 255937 + tpg|BK006942.2| 256024 - INS 
 tpg|BK006942.2| 96077 + tpg|BK006942.2| 95611 - INS 
 tpg|BK006942.2| 134637 + tpg|BK006942.2| 134554 - INS 
 tpg|BK006942.2| 432544 + tpg|BK006942.2| 431886 - INS 
 tpg|BK006942.2| 243246 + tpg|BK006942.2| 243073 - INS 
 tpg|BK006942.2| 363947 + tpg|BK006942.2| 363524 - INS 
 tpg|BK006942.2| 83162 + tpg|BK006942.2| 82703 - INS 
 tpg|BK006942.2| 29771 + tpg|BK006942.2| 29590 - INS 
 tpg|BK006942.2| 26520 + tpg|BK006942.2| 26250 - INS 
 tpg|BK006942.2| 25315 + tpg|BK006942.2| 24952 - INS 
 tpg|BK006942.2| 170949 + tpg|BK006942.2| 171633 - INS 
 tpg|BK006942.2| 145103 + tpg|BK006942.2| 144347 - INS 
 tpg|BK006942.2| 138179 + tpg|BK006942.2| 137719 - INS 
 tpg|BK006942.2| 286780 + tpg|BK006942.2| 286473 - INS 
 tpg|BK006942.2| 119166 + tpg|BK006942.2| 118665 - INS 
 tpg|BK006942.2| 190544 + tpg|BK006942.2| 190136 - INS 
 tpg|BK006942.2| 102233 + tpg|BK006942.2| 101998 - INS 
 tpg|BK006942.2| 193551 + tpg|BK006942.2| 193659 - INS 
 tpg|BK006942.2| 264941 + tpg|BK006942.2| 264779 - INS 
 tpg|BK006942.2| 99374 + tpg|BK006942.2| 99412 - INS 
 tpg|BK006942.2| 314174 + tpg|BK006942.2| 314111 - INS 
 tpg|BK006942.2| 86742 + tpg|BK006942.2| 86399 - INS 
 tpg|BK006942.2| 262936 + tpg|BK006942.2| 262900 - INS 
 tpg|BK006942.2| 57896 + tpg|BK006942.2| 57657 - INS 
 tpg|BK006942.2| 269640 + tpg|BK006942.2| 269425 - INS 
 tpg|BK006942.2| 185729 + tpg|BK006942.2| 185252 - INS 
 tpg|BK006942.2| 192738 + tpg|BK006942.2| 192072 - INS 
 tpg|BK006942.2| 89620 + tpg|BK006942.2| 89286 - INS 
 tpg|BK006942.2| 173198 + tpg|BK006942.2| 172942 - INS 
 tpg|BK006942.2| 355088 + tpg|BK006942.2| 354597 - INS 
 tpg|BK006942.2| 436713 + tpg|BK006942.2| 436114 - INS 
 tpg|BK006942.2| 329390 + tpg|BK006942.2| 329183 - INS 
 tpg|BK006942.2| 358229 + tpg|BK006942.2| 358605 - INS 
 tpg|BK006942.2| 375409 + tpg|BK006942.2| 375283 - INS 
 tpg|BK006942.2| 34023 + tpg|BK006942.2| 33455 - INS 
 tpg|BK006942.2| 20420 + tpg|BK006942.2| 20300 - INS 
 tpg|BK006942.2| 129976 + tpg|BK006942.2| 129377 - INS 
 tpg|BK006942.2| 426094 + tpg|BK006942.2| 425524 - INS 
 tpg|BK006942.2| 27603 + tpg|BK006942.2| 28157 - INS 
 tpg|BK006942.2| 418421 + tpg|BK006942.2| 418615 - INS 
 tpg|BK006942.2| 34545 + tpg|BK006942.2| 35076 - INS 
 tpg|BK006942.2| 292161 + tpg|BK006942.2| 291846 - INS 
 tpg|BK006942.2| 174071 + tpg|BK006942.2| 173531 - INS 
 tpg|BK006942.2| 275513 + tpg|BK006942.2| 275599 - INS 
 tpg|BK006942.2| 185103 + tpg|BK006942.2| 184742 - INS 
 tpg|BK006942.2| 186608 + tpg|BK006942.2| 186623 - INS 
 tpg|BK006942.2| 110531 + tpg|BK006942.2| 110279 - INS 
 tpg|BK006942.2| 238224 + tpg|BK006942.2| 238118 - INS 
 tpg|BK006942.2| 377877 + tpg|BK006942.2| 377512 - INS 
 tpg|BK006942.2| 324129 + tpg|BK006942.2| 324757 - INS 
 tpg|BK006942.2| 295811 + tpg|BK006942.2| 296410 - INS 
 tpg|BK006942.2| 24445 + tpg|BK006942.2| 23912 - INS 
 tpg|BK006942.2| 345978 + tpg|BK006942.2| 345681 - INS 
 tpg|BK006942.2| 350866 + tpg|BK006942.2| 350766 - INS 
 tpg|BK006942.2| 336435 + tpg|BK006942.2| 336110 - INS 
 tpg|BK006942.2| 142269 + tpg|BK006942.2| 142000 - INS 
 tpg|BK006942.2| 38347 + tpg|BK006942.2| 38093 - INS 
 tpg|BK006942.2| 407307 + tpg|BK006942.2| 406954 - INS 
 tpg|BK006942.2| 367691 + tpg|BK006942.2| 368146 - INS 
 tpg|BK006942.2| 107877 + tpg|BK006942.2| 108359 - INS 
 tpg|BK006942.2| 348660 + tpg|BK006942.2| 348241 - INS 
 tpg|BK006942.2| 436004 + tpg|BK006942.2| 435338 - INS 
 tpg|BK006942.2| 293871 + tpg|BK006942.2| 294098 - INS 
 tpg|BK006942.2| 338271 + tpg|BK006942.2| 338053 - INS 
 tpg|BK006942.2| 95197 + tpg|BK006942.2| 95051 - INS 
 tpg|BK006942.2| 309082 + tpg|BK006942.2| 308497 - INS 
 tpg|BK006942.2| 181732 + tpg|BK006942.2| 181494 - INS 
 tpg|BK006942.2| 124362 + tpg|BK006942.2| 123898 - INS 
 tpg|BK006942.2| 92049 + tpg|BK006942.2| 91335 - INS 
 tpg|BK006942.2| 381584 + tpg|BK006942.2| 381281 - INS 
 tpg|BK006942.2| 65531 + tpg|BK006942.2| 65232 - INS 
 tpg|BK006942.2| 174573 + tpg|BK006942.2| 174444 - INS 
 tpg|BK006942.2| 42854 + tpg|BK006942.2| 42143 - INS 
 tpg|BK006942.2| 363067 + tpg|BK006942.2| 363115 - INS 
 tpg|BK006942.2| 170229 + tpg|BK006942.2| 170636 - INS 
 tpg|BK006942.2| 68137 + tpg|BK006942.2| 67960 - INS 
 tpg|BK006942.2| 346611 + tpg|BK006942.2| 346887 - INS 
 tpg|BK006942.2| 209655 + tpg|BK006942.2| 209275 - INS 
 tpg|BK006942.2| 182258 + tpg|BK006942.2| 182662 - INS 
 tpg|BK006942.2| 66324 + tpg|BK006942.2| 66105 - INS 
 tpg|BK006942.2| 208405 + tpg|BK006942.2| 208190 - INS 
 tpg|BK006942.2| 219241 + tpg|BK006942.2| 218749 - INS 
 tpg|BK006942.2| 119781 + tpg|BK006942.2| 120086 - INS 
 tpg|BK006942.2| 260169 + tpg|BK006942.2| 260035 - INS 
 tpg|BK006942.2| 372209 + tpg|BK006942.2| 372039 - INS 
 tpg|BK006942.2| 38982 + tpg|BK006942.2| 38769 - INS 
 tpg|BK006942.2| 226826 + tpg|BK006942.2| 226533 - INS TA
 tpg|BK006935.2| 76987 + tpg|BK006935.2| 77541 - INS 
 tpg|BK006935.2| 191422 + tpg|BK006935.2| 191037 - INS 
 tpg|BK006935.2| 33474 + tpg|BK006935.2| 33724 - INS 
 tpg|BK006935.2| 148636 + tpg|BK006935.2| 148268 - INS 
 tpg|BK006935.2| 37093 + tpg|BK006935.2| 37226 - INS 
 tpg|BK006935.2| 82441 + tpg|BK006935.2| 83091 - INS 
 tpg|BK006935.2| 125576 + tpg|BK006935.2| 126075 - INS 
 tpg|BK006935.2| 74918 + tpg|BK006935.2| 75613 - INS 
 tpg|BK006937.2| 50606 + tpg|BK006937.2| 50957 - INS 
 tpg|BK006935.2| 193066 + tpg|BK006935.2| 192538 - INS 
 tpg|BK006935.2| 13009 + tpg|BK006935.2| 12886 - INS 
 tpg|BK006935.2| 40668 + tpg|BK006935.2| 40356 - INS 
 tpg|BK006935.2| 195793 + tpg|BK006935.2| 195703 - INS 
 tpg|BK006935.2| 53168 + tpg|BK006935.2| 53466 - INS 
 tpg|BK006935.2| 57652 + tpg|BK006935.2| 58052 - INS 
 tpg|BK006935.2| 41904 + tpg|BK006935.2| 41316 - INS 
 tpg|BK006935.2| 116599 + tpg|BK006935.2| 116236 - INS 
 tpg|BK006935.2| 186416 + tpg|BK006935.2| 187137 - INS 
 tpg|BK006935.2| 228932 + tpg|BK006935.2| 229096 - INS 
 tpg|BK006935.2| 113525 + tpg|BK006935.2| 113017 - INS 
 tpg|BK006935.2| 156990 + tpg|BK006935.2| 156403 - INS 
 tpg|BK006935.2| 115153 + tpg|BK006935.2| 114617 - INS 
 tpg|BK006935.2| 110669 + tpg|BK006935.2| 110649 - INS 
 tpg|BK006935.2| 227524 + tpg|BK006935.2| 227819 - INS 
 tpg|BK006935.2| 72985 + tpg|BK006935.2| 73627 - INS 
 tpg|BK006935.2| 109751 + tpg|BK006935.2| 109413 - INS 
 tpg|BK006935.2| 1553 + tpg|BK006935.2| 1707 - INS 
 tpg|BK006935.2| 131264 + tpg|BK006935.2| 130988 - INS 
 tpg|BK006935.2| 66219 + tpg|BK006935.2| 66836 - INS 
 tpg|BK006935.2| 31851 + tpg|BK006935.2| 32059 - INS 
 tpg|BK006935.2| 127092 + tpg|BK006935.2| 126961 - INS 
 tpg|BK006935.2| 96428 + tpg|BK006935.2| 96106 - INS 
 tpg|BK006935.2| 49972 + tpg|BK006935.2| 49957 - INS 
 tpg|BK006935.2| 35924 + tpg|BK006935.2| 36605 - INS 
 tpg|BK006935.2| 86472 + tpg|BK006935.2| 86892 - INS 
 tpg|BK006935.2| 119369 + tpg|BK006935.2| 119504 - INS 
 tpg|BK006935.2| 10080 + tpg|BK006935.2| 9458 - INS 
 tpg|BK006935.2| 61189 + tpg|BK006935.2| 60683 - INS 
 tpg|BK006935.2| 65304 + tpg|BK006935.2| 65938 - INS 
 tpg|BK006935.2| 68990 + tpg|BK006935.2| 68404 - INS 
 tpg|BK006935.2| 136676 + tpg|BK006935.2| 136554 - INS 
 tpg|BK006935.2| 107692 + tpg|BK006935.2| 107313 - INS 
 tpg|BK006935.2| 60152 + tpg|BK006935.2| 60042 - INS 
 tpg|BK006935.2| 130047 + tpg|BK006935.2| 129517 - INS 
 tpg|BK006935.2| 170234 + tpg|BK006935.2| 169653 - INS 
 tpg|BK006935.2| 81112 + tpg|BK006935.2| 80567 - INS 
 tpg|BK006935.2| 198413 + tpg|BK006935.2| 198891 - INS 
 tpg|BK006935.2| 180279 + tpg|BK006935.2| 179944 - INS 
 tpg|BK006935.2| 132051 + tpg|BK006935.2| 132067 - INS 
 tpg|BK006935.2| 133409 + tpg|BK006935.2| 133062 - INS 
 tpg|BK006935.2| 171875 + tpg|BK006935.2| 171296 - INS 
 tpg|BK006935.2| 150394 + tpg|BK006935.2| 149647 - INS 
 tpg|BK006935.2| 44465 + tpg|BK006935.2| 44240 - INS 
 tpg|BK006935.2| 99216 + tpg|BK006935.2| 98558 - INS 
 tpg|BK006935.2| 124719 + tpg|BK006935.2| 124133 - INS 
 tpg|BK006935.2| 52360 + tpg|BK006935.2| 51711 - INS 
 tpg|BK006935.2| 7024 + tpg|BK006935.2| 6934 - INS 
 tpg|BK006935.2| 38761 + tpg|BK006935.2| 38266 - INS 
 tpg|BK006935.2| 16847 + tpg|BK006935.2| 16576 - INS 
 tpg|BK006935.2| 102461 + tpg|BK006935.2| 102303 - INS 
 tpg|BK006935.2| 155669 + tpg|BK006935.2| 154897 - INS 
 tpg|BK006935.2| 175140 + tpg|BK006935.2| 175213 - INS 
 tpg|BK006935.2| 95287 + tpg|BK006935.2| 95344 - INS 
 tpg|BK006935.2| 177214 + tpg|BK006935.2| 176709 - INS 
 tpg|BK006935.2| 35406 + tpg|BK006935.2| 35073 - INS 
 tpg|BK006935.2| 184358 + tpg|BK006935.2| 184097 - INS 
 tpg|BK006935.2| 134474 + tpg|BK006935.2| 134375 - INS 
 tpg|BK006935.2| 167490 + tpg|BK006935.2| 166827 - INS 
 tpg|BK006935.2| 8535 + tpg|BK006935.2| 8638 - INS 
 tpg|BK006935.2| 153275 + tpg|BK006935.2| 152724 - INS 
 tpg|BK006935.2| 72159 + tpg|BK006935.2| 72044 - INS 
 tpg|BK006935.2| 141727 + tpg|BK006935.2| 141223 - INS 
 tpg|BK006935.2| 7715 + tpg|BK006935.2| 7417 - INS 
 tpg|BK006935.2| 21625 + tpg|BK006935.2| 21319 - INS 
 tpg|BK006935.2| 20823 + tpg|BK006935.2| 20751 - INS 
 tpg|BK006935.2| 88096 + tpg|BK006935.2| 87415 - INS 
 tpg|BK006935.2| 122646 + tpg|BK006935.2| 122502 - INS 
 tpg|BK006935.2| 42847 + tpg|BK006935.2| 43151 - INS 
 tpg|BK006935.2| 112036 + tpg|BK006935.2| 111785 - INS 
 tpg|BK006935.2| 19000 + tpg|BK006935.2| 18841 - INS 
 tpg|BK006935.2| 142322 + tpg|BK006935.2| 142020 - INS 
 tpg|BK006935.2| 151326 + tpg|BK006935.2| 151121 - INS 
 tpg|BK006935.2| 137925 + tpg|BK006935.2| 137294 - INS 
 tpg|BK006935.2| 63401 + tpg|BK006935.2| 63026 - INS 
 tpg|BK006935.2| 196817 + tpg|BK006935.2| 196488 - INS 
 tpg|BK006935.2| 90952 + tpg|BK006935.2| 90904 - INS 
 tpg|BK006935.2| 177564 + tpg|BK006935.2| 177874 - INS 
 tpg|BK006935.2| 179013 + tpg|BK006935.2| 178887 - INS 
 tpg|BK006935.2| 48692 + tpg|BK006935.2| 48354 - INS 
 tpg|BK006935.2| 69770 + tpg|BK006935.2| 69620 - INS 
 tpg|BK006935.2| 56293 + tpg|BK006935.2| 55952 - INS 
 tpg|BK006935.2| 185447 + tpg|BK006935.2| 185165 - INS 
 tpg|BK006935.2| 121179 + tpg|BK006935.2| 120712 - INS 
 tpg|BK006935.2| 168841 + tpg|BK006935.2| 168651 - INS 
 tpg|BK006935.2| 47849 + tpg|BK006935.2| 47186 - INS 
 tpg|BK006935.2| 92370 + tpg|BK006935.2| 92188 - INS 
 tpg|BK006935.2| 144004 + tpg|BK006935.2| 143299 - INS 
 tpg|BK006935.2| 138502 + tpg|BK006935.2| 138366 - INS 
 tpg|BK006935.2| 174220 + tpg|BK006935.2| 173653 - INS 
 tpg|BK006935.2| 153664 + tpg|BK006935.2| 153299 - INS 
 tpg|BK006935.2| 99843 + tpg|BK006935.2| 99525 - INS 
 tpg|BK006935.2| 207805 + tpg|BK006935.2| 207320 - INS TACG
 tpg|BK006935.2| 94060 + tpg|BK006935.2| 93672 - INS 
 tpg|BK006935.2| 93147 + tpg|BK006935.2| 92747 - INS 
 tpg|BK006935.2| 85874 + tpg|BK006935.2| 85395 - INS 
 tpg|BK006935.2| 84725 + tpg|BK006935.2| 84542 - INS 
 tpg|BK006935.2| 56877 + tpg|BK006935.2| 56618 - INS 
 tpg|BK006935.2| 193411 + tpg|BK006935.2| 193686 - INS 
 tpg|BK006935.2| 200217 + tpg|BK006935.2| 200763 - INS 
 tpg|BK006935.2| 64695 + tpg|BK006935.2| 64199 - INS 
 tpg|BK006935.2| 78857 + tpg|BK006935.2| 78095 - INS 
 tpg|BK006935.2| 209009 + tpg|BK006935.2| 209601 - INS 
 tpg|BK006935.2| 128078 + tpg|BK006935.2| 128836 - INS 
 tpg|BK006935.2| 189911 + tpg|BK006935.2| 190159 - INS 
 tpg|BK006935.2| 145786 + tpg|BK006935.2| 145880 - INS 
 tpg|BK006935.2| 201946 + tpg|BK006935.2| 201243 - INS 
 tpg|BK006935.2| 11012 + tpg|BK006935.2| 11259 - INS 
 tpg|BK006935.2| 29749 + tpg|BK006935.2| 30503 - INS 
 tpg|BK006935.2| 188130 + tpg|BK006935.2| 187650 - INS 
 tpg|BK006935.2| 13702 + tpg|BK006935.2| 14024 - INS 
 tpg|BK006935.2| 177963 + tpg|BK006935.2| 178521 - INS 
 tpg|BK006935.2| 130465 + tpg|BK006935.2| 130358 - INS 
 tpg|BK006935.2| 79483 + tpg|BK006935.2| 79311 - INS 
 tpg|BK006935.2| 89983 + tpg|BK006935.2| 90360 - INS 
 tpg|BK006935.2| 168120 + tpg|BK006935.2| 167849 - INS 
 tpg|BK006935.2| 70809 + tpg|BK006935.2| 70531 - INS 
 tpg|BK006937.2| 59352 + tpg|BK006937.2| 58845 - INS 
 tpg|BK006937.2| 122408 + tpg|BK006937.2| 122192 - INS 
 tpg|BK006937.2| 270542 + tpg|BK006937.2| 270799 - INS 
 tpg|BK006937.2| 224465 + tpg|BK006937.2| 224780 - INS 
 tpg|BK006937.2| 1914 + tpg|BK006937.2| 1997 - INS 
 tpg|BK006937.2| 63481 + tpg|BK006937.2| 63327 - INS 
 tpg|BK006937.2| 229628 + tpg|BK006937.2| 228973 - INS 
 tpg|BK006937.2| 198721 + tpg|BK006937.2| 197961 - INS 
 tpg|BK006937.2| 209176 + tpg|BK006937.2| 209781 - INS 
 tpg|BK006937.2| 210859 + tpg|BK006937.2| 210829 - INS 
 tpg|BK006937.2| 94243 + tpg|BK006937.2| 93883 - INS 
 tpg|BK006937.2| 106860 + tpg|BK006937.2| 106965 - INS 
 tpg|BK006937.2| 152910 + tpg|BK006937.2| 153240 - INS 
 tpg|BK006937.2| 267645 + tpg|BK006937.2| 267683 - INS 
 tpg|BK006937.2| 282074 + tpg|BK006937.2| 282022 - INS 
 tpg|BK006937.2| 247761 + tpg|BK006937.2| 247348 - INS 
 tpg|BK006937.2| 178133 + tpg|BK006937.2| 178627 - INS 
 tpg|BK006937.2| 67639 + tpg|BK006937.2| 67698 - INS 
 tpg|BK006937.2| 271787 + tpg|BK006937.2| 271445 - INS 
 tpg|BK006937.2| 47480 + tpg|BK006937.2| 47006 - INS 
 tpg|BK006937.2| 234598 + tpg|BK006937.2| 234415 - INS 
 tpg|BK006937.2| 57251 + tpg|BK006937.2| 57886 - INS 
 tpg|BK006937.2| 918 + tpg|BK006937.2| 715 - INS 
 tpg|BK006937.2| 175384 + tpg|BK006937.2| 175192 - INS 
 tpg|BK006937.2| 41300 + tpg|BK006937.2| 40525 - INS 
 tpg|BK006937.2| 225903 + tpg|BK006937.2| 225173 - INS 
 tpg|BK006937.2| 73432 + tpg|BK006937.2| 73301 - INS 
 tpg|BK006937.2| 35004 + tpg|BK006937.2| 35674 - INS 
 tpg|BK006934.2| 58433 + tpg|BK006934.2| 58966 - INS 
 tpg|BK006937.2| 239948 + tpg|BK006937.2| 239924 - INS 
 tpg|BK006934.2| 49785 + tpg|BK006934.2| 49555 - INS 
 tpg|BK006937.2| 264898 + tpg|BK006937.2| 264132 - INS 
 tpg|BK006937.2| 288031 + tpg|BK006937.2| 287825 - INS 
 tpg|BK006934.2| 490415 + tpg|BK006934.2| 490928 - INS 
 tpg|BK006937.2| 70790 + tpg|BK006937.2| 70026 - INS 
 tpg|BK006934.2| 69809 + tpg|BK006934.2| 70224 - INS 
 tpg|BK006937.2| 166465 + tpg|BK006937.2| 165706 - INS 
 tpg|BK006937.2| 55977 + tpg|BK006937.2| 56341 - INS 
 tpg|BK006934.2| 482357 + tpg|BK006934.2| 481725 - INS 
 tpg|BK006937.2| 54127 + tpg|BK006937.2| 53428 - INS 
 tpg|BK006934.2| 366038 + tpg|BK006934.2| 366642 - INS 
 tpg|BK006937.2| 206631 + tpg|BK006937.2| 206834 - INS 
 tpg|BK006934.2| 175225 + tpg|BK006934.2| 174968 - INS 
 tpg|BK006937.2| 296919 + tpg|BK006937.2| 297191 - INS 
 tpg|BK006934.2| 242947 + tpg|BK006934.2| 243714 - INS 
 tpg|BK006937.2| 279372 + tpg|BK006937.2| 278981 - INS 
 tpg|BK006937.2| 295915 + tpg|BK006937.2| 295340 - INS 
 tpg|BK006934.2| 411726 + tpg|BK006934.2| 412280 - INS 
 tpg|BK006937.2| 253583 + tpg|BK006937.2| 253311 - INS 
 tpg|BK006937.2| 309555 + tpg|BK006937.2| 309132 - INS 
 tpg|BK006934.2| 140926 + tpg|BK006934.2| 141622 - INS 
 tpg|BK006934.2| 236850 + tpg|BK006934.2| 237512 - INS 
 tpg|BK006937.2| 241173 + tpg|BK006937.2| 241054 - INS 
 tpg|BK006934.2| 230432 + tpg|BK006934.2| 230016 - INS 
 tpg|BK006937.2| 103503 + tpg|BK006937.2| 103393 - INS 
 tpg|BK006937.2| 101527 + tpg|BK006937.2| 102295 - INS 
 tpg|BK006934.2| 477926 + tpg|BK006934.2| 477560 - INS 
 tpg|BK006937.2| 97656 + tpg|BK006937.2| 97935 - INS 
 tpg|BK006937.2| 304295 + tpg|BK006937.2| 304320 - INS 
 tpg|BK006934.2| 443827 + tpg|BK006934.2| 444143 - INS 
 tpg|BK006937.2| 233309 + tpg|BK006937.2| 233727 - INS 
 tpg|BK006934.2| 176622 + tpg|BK006934.2| 177035 - INS 
 tpg|BK006937.2| 81379 + tpg|BK006937.2| 80811 - INS 
 tpg|BK006934.2| 160044 + tpg|BK006934.2| 159686 - INS 
 tpg|BK006937.2| 274260 + tpg|BK006937.2| 273950 - INS 
 tpg|BK006934.2| 482777 + tpg|BK006934.2| 482299 - INS 
 tpg|BK006937.2| 312532 + tpg|BK006937.2| 313009 - INS 
 tpg|BK006937.2| 154634 + tpg|BK006937.2| 154190 - INS 
 tpg|BK006934.2| 98594 + tpg|BK006934.2| 98291 - INS 
 tpg|BK006937.2| 164785 + tpg|BK006937.2| 165162 - INS 
 tpg|BK006937.2| 15883 + tpg|BK006937.2| 16212 - INS 
 tpg|BK006934.2| 217983 + tpg|BK006934.2| 217971 - INS 
 tpg|BK006937.2| 61999 + tpg|BK006937.2| 61537 - INS 
 tpg|BK006937.2| 211679 + tpg|BK006937.2| 211729 - INS 
 tpg|BK006934.2| 191599 + tpg|BK006934.2| 191672 - INS 
 tpg|BK006937.2| 134626 + tpg|BK006937.2| 134682 - INS 
 tpg|BK006937.2| 44522 + tpg|BK006937.2| 44167 - INS 
 tpg|BK006934.2| 196790 + tpg|BK006934.2| 196438 - INS 
 tpg|BK006937.2| 106049 + tpg|BK006937.2| 105675 - INS 
 tpg|BK006934.2| 160709 + tpg|BK006934.2| 160381 - INS 
 tpg|BK006937.2| 243387 + tpg|BK006937.2| 242981 - INS 
 tpg|BK006937.2| 61442 + tpg|BK006937.2| 61008 - INS 
 tpg|BK006934.2| 337942 + tpg|BK006934.2| 338187 - INS 
 tpg|BK006937.2| 195553 + tpg|BK006937.2| 195061 - INS 
 tpg|BK006937.2| 230658 + tpg|BK006937.2| 231039 - INS 
 tpg|BK006934.2| 410102 + tpg|BK006934.2| 409958 - INS 
 tpg|BK006937.2| 66332 + tpg|BK006937.2| 66535 - INS 
 tpg|BK006937.2| 167340 + tpg|BK006937.2| 168043 - INS 
 tpg|BK006937.2| 215838 + tpg|BK006937.2| 215627 - INS 
 tpg|BK006937.2| 41801 + tpg|BK006937.2| 41458 - INS 
 tpg|BK006937.2| 236798 + tpg|BK006937.2| 236288 - INS 
 tpg|BK006937.2| 22077 + tpg|BK006937.2| 21731 - INS 
 tpg|BK006937.2| 52283 + tpg|BK006937.2| 52012 - INS 
 tpg|BK006937.2| 238092 + tpg|BK006937.2| 237874 - INS 
 tpg|BK006937.2| 147053 + tpg|BK006937.2| 147607 - INS 
 tpg|BK006937.2| 71282 + tpg|BK006937.2| 71480 - INS 
 tpg|BK006937.2| 288785 + tpg|BK006937.2| 289125 - INS 
 tpg|BK006937.2| 187207 + tpg|BK006937.2| 187826 - INS 
 tpg|BK006937.2| 196231 + tpg|BK006937.2| 195917 - INS 
 tpg|BK006937.2| 14838 + tpg|BK006937.2| 14815 - INS 
 tpg|BK006937.2| 121072 + tpg|BK006937.2| 120800 - INS 
 tpg|BK006937.2| 290332 + tpg|BK006937.2| 289663 - INS 
 tpg|BK006937.2| 45737 + tpg|BK006937.2| 45900 - INS 
 tpg|BK006937.2| 284081 + tpg|BK006937.2| 283855 - INS 
 tpg|BK006937.2| 155035 + tpg|BK006937.2| 155798 - INS 
 tpg|BK006937.2| 189015 + tpg|BK006937.2| 189631 - INS 
 tpg|BK006934.2| 334861 + tpg|BK006934.2| 334773 - INS 
 tpg|BK006934.2| 315989 + tpg|BK006934.2| 315848 - INS 
 tpg|BK006937.2| 17785 + tpg|BK006937.2| 17755 - INS 
 tpg|BK006934.2| 377860 + tpg|BK006934.2| 377760 - INS 
 tpg|BK006937.2| 157693 + tpg|BK006937.2| 157424 - INS 
 tpg|BK006937.2| 172529 + tpg|BK006937.2| 172952 - INS 
 tpg|BK006934.2| 379908 + tpg|BK006934.2| 379235 - INS 
 tpg|BK006937.2| 127145 + tpg|BK006937.2| 126723 - INS 
 tpg|BK006937.2| 216989 + tpg|BK006937.2| 217043 - INS 
 tpg|BK006934.2| 93118 + tpg|BK006934.2| 92530 - INS 
 tpg|BK006937.2| 120072 + tpg|BK006937.2| 119939 - INS 
 tpg|BK006937.2| 94881 + tpg|BK006937.2| 94510 - INS 
 tpg|BK006937.2| 218967 + tpg|BK006937.2| 218892 - INS 
 tpg|BK006937.2| 137697 + tpg|BK006937.2| 137723 - INS 
 tpg|BK006937.2| 104892 + tpg|BK006937.2| 104894 - INS 
 tpg|BK006934.2| 347014 + tpg|BK006934.2| 346776 - INS 
 tpg|BK006937.2| 226757 + tpg|BK006937.2| 226432 - INS 
 tpg|BK006937.2| 37620 + tpg|BK006937.2| 36953 - INS 
 tpg|BK006937.2| 99803 + tpg|BK006937.2| 100473 - INS 
 tpg|BK006934.2| 131037 + tpg|BK006934.2| 130941 - INS 
 tpg|BK006934.2| 463794 + tpg|BK006934.2| 463872 - INS 
 tpg|BK006937.2| 180289 + tpg|BK006937.2| 180019 - INS 
 tpg|BK006937.2| 54936 + tpg|BK006937.2| 55329 - INS 
 tpg|BK006937.2| 48330 + tpg|BK006937.2| 48166 - INS 
 tpg|BK006937.2| 202902 + tpg|BK006937.2| 202760 - INS 
 tpg|BK006937.2| 220808 + tpg|BK006937.2| 220962 - INS 
 tpg|BK006937.2| 82055 + tpg|BK006937.2| 81383 - INS 
 tpg|BK006934.2| 298795 + tpg|BK006934.2| 298411 - INS 
 tpg|BK006937.2| 206038 + tpg|BK006937.2| 205716 - INS 
 tpg|BK006934.2| 38127 + tpg|BK006934.2| 37555 - INS 
 tpg|BK006934.2| 325248 + tpg|BK006934.2| 325911 - INS 
 tpg|BK006937.2| 292121 + tpg|BK006937.2| 291813 - INS 
 tpg|BK006934.2| 263215 + tpg|BK006934.2| 263554 - INS 
 tpg|BK006937.2| 49159 + tpg|BK006937.2| 49559 - INS 
 tpg|BK006934.2| 485788 + tpg|BK006934.2| 486447 - INS 
 tpg|BK006937.2| 24312 + tpg|BK006937.2| 24491 - INS 
 tpg|BK006934.2| 505251 + tpg|BK006934.2| 505583 - INS 
 tpg|BK006937.2| 254181 + tpg|BK006937.2| 254723 - INS 
 tpg|BK006934.2| 120679 + tpg|BK006934.2| 120052 - INS 
 tpg|BK006937.2| 75102 + tpg|BK006937.2| 74407 - INS 
 tpg|BK006937.2| 241838 + tpg|BK006937.2| 241543 - INS 
 tpg|BK006937.2| 277854 + tpg|BK006937.2| 277569 - INS 
 tpg|BK006937.2| 184860 + tpg|BK006937.2| 185380 - INS 
 tpg|BK006934.2| 60068 + tpg|BK006934.2| 59895 - INS 
 tpg|BK006937.2| 129861 + tpg|BK006937.2| 129613 - INS 
 tpg|BK006937.2| 32931 + tpg|BK006937.2| 32905 - INS 
 tpg|BK006934.2| 470218 + tpg|BK006934.2| 470101 - INS 
 tpg|BK006934.2| 507756 + tpg|BK006934.2| 507040 - INS 
 tpg|BK006937.2| 223166 + tpg|BK006937.2| 223057 - INS 
 tpg|BK006937.2| 136069 + tpg|BK006937.2| 135585 - INS 
 tpg|BK006937.2| 249188 + tpg|BK006937.2| 249083 - INS 
 tpg|BK006934.2| 68545 + tpg|BK006934.2| 68784 - INS 
 tpg|BK006937.2| 176701 + tpg|BK006937.2| 176082 - INS 
 tpg|BK006934.2| 279795 + tpg|BK006934.2| 280107 - INS 
 tpg|BK006937.2| 227446 + tpg|BK006937.2| 227275 - INS 
 tpg|BK006937.2| 118514 + tpg|BK006937.2| 118780 - INS 
 tpg|BK006934.2| 272035 + tpg|BK006934.2| 272383 - INS 
 tpg|BK006937.2| 244669 + tpg|BK006937.2| 244529 - INS 
 tpg|BK006937.2| 249626 + tpg|BK006937.2| 249981 - INS 
 tpg|BK006934.2| 461655 + tpg|BK006934.2| 461563 - INS 
 tpg|BK006937.2| 79952 + tpg|BK006937.2| 79686 - INS 
 tpg|BK006937.2| 252035 + tpg|BK006937.2| 251928 - INS 
 tpg|BK006937.2| 266823 + tpg|BK006937.2| 266909 - INS 
 tpg|BK006937.2| 305750 + tpg|BK006937.2| 305198 - INS 
 tpg|BK006934.2| 264086 + tpg|BK006934.2| 264858 - INS TTCATAT
 tpg|BK006937.2| 192495 + tpg|BK006937.2| 192260 - INS 
 tpg|BK006937.2| 11460 + tpg|BK006937.2| 11046 - INS 
 tpg|BK006934.2| 181003 + tpg|BK006934.2| 180667 - INS 
 tpg|BK006934.2| 483477 + tpg|BK006934.2| 483166 - INS 
 tpg|BK006934.2| 221808 + tpg|BK006934.2| 221504 - INS 
 tpg|BK006934.2| 214295 + tpg|BK006934.2| 214209 - INS 
 tpg|BK006934.2| 164567 + tpg|BK006934.2| 164597 - INS 
 tpg|BK006937.2| 310768 + tpg|BK006937.2| 311198 - INS 
 tpg|BK006934.2| 19697 + tpg|BK006934.2| 19212 - INS 
 tpg|BK006937.2| 145352 + tpg|BK006937.2| 144751 - INS 
 tpg|BK006937.2| 286054 + tpg|BK006937.2| 286333 - INS 
 tpg|BK006937.2| 222201 + tpg|BK006937.2| 221479 - INS 
 tpg|BK006934.2| 354144 + tpg|BK006934.2| 354128 - INS 
 tpg|BK006937.2| 108659 + tpg|BK006937.2| 108397 - INS 
 tpg|BK006934.2| 241047 + tpg|BK006934.2| 240757 - INS 
 tpg|BK006937.2| 9413 + tpg|BK006937.2| 9123 - INS 
 tpg|BK006937.2| 286687 + tpg|BK006937.2| 286883 - INS 
 tpg|BK006937.2| 139628 + tpg|BK006937.2| 139578 - INS 
 tpg|BK006937.2| 306578 + tpg|BK006937.2| 305908 - INS 
 tpg|BK006937.2| 245915 + tpg|BK006937.2| 245271 - INS 
 tpg|BK006934.2| 188729 + tpg|BK006934.2| 188829 - INS 
 tpg|BK006937.2| 259052 + tpg|BK006937.2| 259065 - INS 
 tpg|BK006934.2| 162709 + tpg|BK006934.2| 162665 - INS 
 tpg|BK006934.2| 79061 + tpg|BK006934.2| 78778 - INS 
 tpg|BK006937.2| 45192 + tpg|BK006937.2| 44874 - INS 
 tpg|BK006937.2| 30121 + tpg|BK006937.2| 30385 - INS 
 tpg|BK006934.2| 33998 + tpg|BK006934.2| 33904 - INS 
 tpg|BK006937.2| 273460 + tpg|BK006937.2| 273118 - INS 
 tpg|BK006934.2| 313371 + tpg|BK006934.2| 314087 - INS 
 tpg|BK006937.2| 44073 + tpg|BK006937.2| 43462 - INS 
 tpg|BK006937.2| 280529 + tpg|BK006937.2| 280639 - INS 
 tpg|BK006937.2| 68819 + tpg|BK006937.2| 68993 - INS 
 tpg|BK006937.2| 191133 + tpg|BK006937.2| 190884 - INS 
 tpg|BK006934.2| 446959 + tpg|BK006934.2| 446754 - INS 
 tpg|BK006937.2| 257155 + tpg|BK006937.2| 256817 - INS 
 tpg|BK006937.2| 133113 + tpg|BK006937.2| 132660 - INS 
 tpg|BK006937.2| 298467 + tpg|BK006937.2| 298584 - INS 
 tpg|BK006937.2| 140409 + tpg|BK006937.2| 140265 - INS 
 tpg|BK006937.2| 136404 + tpg|BK006937.2| 137007 - INS 
 tpg|BK006937.2| 138567 + tpg|BK006937.2| 138556 - INS 
 tpg|BK006934.2| 153908 + tpg|BK006934.2| 154522 - INS 
 tpg|BK006937.2| 124548 + tpg|BK006937.2| 124447 - INS 
 tpg|BK006934.2| 100389 + tpg|BK006934.2| 99628 - INS 
 tpg|BK006937.2| 223931 + tpg|BK006937.2| 223589 - INS 
 tpg|BK006937.2| 307413 + tpg|BK006937.2| 307755 - INS 
 tpg|BK006934.2| 10290 + tpg|BK006934.2| 10089 - INS 
 tpg|BK006937.2| 114539 + tpg|BK006937.2| 113875 - INS 
 tpg|BK006937.2| 282806 + tpg|BK006937.2| 283003 - INS 
 tpg|BK006934.2| 284318 + tpg|BK006934.2| 284645 - INS 
 tpg|BK006937.2| 95790 + tpg|BK006937.2| 95828 - INS 
 tpg|BK006934.2| 275809 + tpg|BK006934.2| 275449 - INS 
 tpg|BK006937.2| 38433 + tpg|BK006937.2| 37697 - INS 
 tpg|BK006937.2| 162074 + tpg|BK006937.2| 161391 - INS 
 tpg|BK006937.2| 115186 + tpg|BK006937.2| 114748 - INS 
 tpg|BK006934.2| 31452 + tpg|BK006934.2| 31132 - INS 
 tpg|BK006937.2| 300272 + tpg|BK006937.2| 299914 - INS 
 tpg|BK006934.2| 487960 + tpg|BK006934.2| 487698 - INS 
 tpg|BK006937.2| 183035 + tpg|BK006937.2| 183266 - INS 
 tpg|BK006937.2| 193605 + tpg|BK006937.2| 193900 - INS 
 tpg|BK006937.2| 272322 + tpg|BK006937.2| 271978 - INS 
 tpg|BK006934.2| 350410 + tpg|BK006934.2| 350654 - INS 
 tpg|BK006937.2| 109230 + tpg|BK006937.2| 109280 - INS 
 tpg|BK006937.2| 291061 + tpg|BK006937.2| 291192 - INS 
 tpg|BK006934.2| 360286 + tpg|BK006934.2| 361046 - INS 
 tpg|BK006937.2| 142581 + tpg|BK006937.2| 141894 - INS 
 tpg|BK006937.2| 93508 + tpg|BK006937.2| 93404 - INS 
 tpg|BK006937.2| 18817 + tpg|BK006937.2| 18182 - INS 
 tpg|BK006937.2| 23410 + tpg|BK006937.2| 22762 - INS 
 tpg|BK006937.2| 255638 + tpg|BK006937.2| 255545 - INS 
 tpg|BK006937.2| 201895 + tpg|BK006937.2| 202038 - INS 
 tpg|BK006937.2| 31947 + tpg|BK006937.2| 31762 - INS 
 tpg|BK006934.2| 512687 + tpg|BK006934.2| 512662 - INS 
 tpg|BK006937.2| 22587 + tpg|BK006937.2| 22139 - INS 
 tpg|BK006937.2| 31441 + tpg|BK006937.2| 31033 - INS 
 tpg|BK006934.2| 143778 + tpg|BK006934.2| 143911 - INS 
 tpg|BK006937.2| 38801 + tpg|BK006937.2| 38214 - INS 
 tpg|BK006937.2| 188646 + tpg|BK006937.2| 189121 - INS 
 tpg|BK006937.2| 212940 + tpg|BK006937.2| 212654 - INS 
 tpg|BK006937.2| 62406 + tpg|BK006937.2| 62586 - INS 
 tpg|BK006937.2| 262681 + tpg|BK006937.2| 261954 - INS 
 tpg|BK006937.2| 197151 + tpg|BK006937.2| 196857 - INS 
 tpg|BK006937.2| 269764 + tpg|BK006937.2| 269612 - INS 
 tpg|BK006937.2| 292760 + tpg|BK006937.2| 292686 - INS 
 tpg|BK006937.2| 237429 + tpg|BK006937.2| 236893 - INS 
 tpg|BK006937.2| 160144 + tpg|BK006937.2| 160175 - INS 
 tpg|BK006937.2| 222594 + tpg|BK006937.2| 222368 - INS 
 tpg|BK006937.2| 265713 + tpg|BK006937.2| 265430 - INS CTGA
 tpg|BK006937.2| 76929 + tpg|BK006937.2| 76837 - INS 
 tpg|BK006937.2| 299681 + tpg|BK006937.2| 299296 - INS 
 tpg|BK006937.2| 158229 + tpg|BK006937.2| 158648 - INS 
 tpg|BK006937.2| 269196 + tpg|BK006937.2| 268848 - INS 
 tpg|BK006937.2| 117184 + tpg|BK006937.2| 117434 - INS 
 tpg|BK006937.2| 6498 + tpg|BK006937.2| 5989 - INS 
 tpg|BK006937.2| 111722 + tpg|BK006937.2| 111289 - INS 
 tpg|BK006937.2| 75861 + tpg|BK006937.2| 75512 - INS 
 tpg|BK006937.2| 248209 + tpg|BK006937.2| 248613 - INS 
 tpg|BK006937.2| 180823 + tpg|BK006937.2| 180595 - INS 
 tpg|BK006934.2| 459851 + tpg|BK006934.2| 459306 - INS 
 tpg|BK006934.2| 396958 + tpg|BK006934.2| 397521 - INS 
 tpg|BK006934.2| 391626 + tpg|BK006934.2| 391373 - INS 
 tpg|BK006934.2| 222362 + tpg|BK006934.2| 221946 - INS 
 tpg|BK006934.2| 209034 + tpg|BK006934.2| 208905 - INS 
 tpg|BK006934.2| 171735 + tpg|BK006934.2| 171077 - INS 
 tpg|BK006934.2| 266724 + tpg|BK006934.2| 266204 - INS 
 tpg|BK006934.2| 420548 + tpg|BK006934.2| 419998 - INS 
 tpg|BK006934.2| 114774 + tpg|BK006934.2| 115194 - INS 
 tpg|BK006934.2| 452649 + tpg|BK006934.2| 452798 - INS 
 tpg|BK006934.2| 394170 + tpg|BK006934.2| 394300 - INS 
 tpg|BK006934.2| 65251 + tpg|BK006934.2| 64620 - INS 
 tpg|BK006934.2| 307246 + tpg|BK006934.2| 307412 - INS 
 tpg|BK006934.2| 46794 + tpg|BK006934.2| 47419 - INS 
 tpg|BK006934.2| 201563 + tpg|BK006934.2| 200970 - INS 
 tpg|BK006934.2| 145040 + tpg|BK006934.2| 144794 - INS 
 tpg|BK006934.2| 500021 + tpg|BK006934.2| 499298 - INS 
 tpg|BK006934.2| 514244 + tpg|BK006934.2| 513568 - INS 
 tpg|BK006934.2| 51823 + tpg|BK006934.2| 51448 - INS 
 tpg|BK006934.2| 352365 + tpg|BK006934.2| 351608 - INS 
 tpg|BK006934.2| 326875 + tpg|BK006934.2| 326932 - INS 
 tpg|BK006934.2| 501449 + tpg|BK006934.2| 501050 - INS 
 tpg|BK006934.2| 281633 + tpg|BK006934.2| 281647 - INS 
 tpg|BK006934.2| 330398 + tpg|BK006934.2| 330549 - INS 
 tpg|BK006934.2| 205237 + tpg|BK006934.2| 204945 - INS 
 tpg|BK006934.2| 383467 + tpg|BK006934.2| 382831 - INS 
 tpg|BK006934.2| 450654 + tpg|BK006934.2| 450178 - INS 
 tpg|BK006934.2| 152589 + tpg|BK006934.2| 152634 - INS 
 tpg|BK006934.2| 312777 + tpg|BK006934.2| 312054 - INS 
 tpg|BK006934.2| 406746 + tpg|BK006934.2| 406725 - INS 
 tpg|BK006934.2| 113835 + tpg|BK006934.2| 113513 - INS 
 tpg|BK006934.2| 112680 + tpg|BK006934.2| 112797 - INS 
 tpg|BK006934.2| 204205 + tpg|BK006934.2| 204452 - INS 
 tpg|BK006934.2| 189754 + tpg|BK006934.2| 189287 - INS 
 tpg|BK006934.2| 386017 + tpg|BK006934.2| 386178 - INS 
 tpg|BK006934.2| 404975 + tpg|BK006934.2| 404377 - INS 
 tpg|BK006934.2| 519532 + tpg|BK006934.2| 519044 - INS 
 tpg|BK006934.2| 309025 + tpg|BK006934.2| 308763 - INS 
 tpg|BK006934.2| 437338 + tpg|BK006934.2| 436963 - INS 
 tpg|BK006934.2| 37183 + tpg|BK006934.2| 37141 - INS 
 tpg|BK006934.2| 433080 + tpg|BK006934.2| 432729 - INS 
 tpg|BK006934.2| 423673 + tpg|BK006934.2| 423235 - INS 
 tpg|BK006934.2| 395552 + tpg|BK006934.2| 394946 - INS 
 tpg|BK006934.2| 74339 + tpg|BK006934.2| 74214 - INS 
 tpg|BK006934.2| 478914 + tpg|BK006934.2| 478151 - INS 
 tpg|BK006934.2| 40536 + tpg|BK006934.2| 39781 - INS 
 tpg|BK006934.2| 116122 + tpg|BK006934.2| 115831 - INS 
 tpg|BK006934.2| 133661 + tpg|BK006934.2| 134427 - INS 
 tpg|BK006934.2| 418565 + tpg|BK006934.2| 418830 - INS 
 tpg|BK006934.2| 396136 + tpg|BK006934.2| 396095 - INS 
 tpg|BK006934.2| 364026 + tpg|BK006934.2| 363900 - INS 
 tpg|BK006934.2| 356842 + tpg|BK006934.2| 356685 - INS 
 tpg|BK006934.2| 94954 + tpg|BK006934.2| 94400 - INS 
 tpg|BK006934.2| 317438 + tpg|BK006934.2| 317619 - INS 
 tpg|BK006934.2| 73053 + tpg|BK006934.2| 73257 - INS 
 tpg|BK006934.2| 441364 + tpg|BK006934.2| 441418 - INS 
 tpg|BK006934.2| 389171 + tpg|BK006934.2| 389659 - INS 
 tpg|BK006934.2| 14478 + tpg|BK006934.2| 14017 - INS 
 tpg|BK006934.2| 42642 + tpg|BK006934.2| 42265 - INS 
 tpg|BK006934.2| 340395 + tpg|BK006934.2| 339756 - INS 
 tpg|BK006934.2| 472402 + tpg|BK006934.2| 471665 - INS 
 tpg|BK006934.2| 197494 + tpg|BK006934.2| 197449 - INS 
 tpg|BK006934.2| 327710 + tpg|BK006934.2| 328122 - INS 
 tpg|BK006934.2| 516294 + tpg|BK006934.2| 515934 - INS 
 tpg|BK006934.2| 55542 + tpg|BK006934.2| 55858 - INS 
 tpg|BK006934.2| 276601 + tpg|BK006934.2| 277293 - INS 
 tpg|BK006934.2| 300868 + tpg|BK006934.2| 301357 - INS 
 tpg|BK006934.2| 5414 + tpg|BK006934.2| 4801 - INS 
 tpg|BK006934.2| 369756 + tpg|BK006934.2| 369509 - INS 
 tpg|BK006934.2| 249885 + tpg|BK006934.2| 249603 - INS 
 tpg|BK006934.2| 124938 + tpg|BK006934.2| 124804 - INS 
 tpg|BK006934.2| 247288 + tpg|BK006934.2| 247067 - INS 
 tpg|BK006934.2| 402610 + tpg|BK006934.2| 402377 - INS 
 tpg|BK006934.2| 467133 + tpg|BK006934.2| 467267 - INS 
 tpg|BK006934.2| 368186 + tpg|BK006934.2| 368010 - INS 
 tpg|BK006934.2| 118010 + tpg|BK006934.2| 118016 - INS 
 tpg|BK006934.2| 361923 + tpg|BK006934.2| 362550 - INS 
 tpg|BK006934.2| 75610 + tpg|BK006934.2| 74979 - INS 
 tpg|BK006934.2| 321682 + tpg|BK006934.2| 321265 - INS 
 tpg|BK006934.2| 71895 + tpg|BK006934.2| 71567 - INS 
 tpg|BK006934.2| 107410 + tpg|BK006934.2| 107387 - INS 
 tpg|BK006934.2| 208249 + tpg|BK006934.2| 207862 - INS 
 tpg|BK006934.2| 341733 + tpg|BK006934.2| 341670 - INS 
 tpg|BK006934.2| 415673 + tpg|BK006934.2| 415735 - INS 
 tpg|BK006934.2| 382407 + tpg|BK006934.2| 381801 - INS 
 tpg|BK006934.2| 262340 + tpg|BK006934.2| 262756 - INS 
 tpg|BK006934.2| 399089 + tpg|BK006934.2| 399304 - INS 
 tpg|BK006934.2| 32016 + tpg|BK006934.2| 31873 - INS 
 tpg|BK006934.2| 302513 + tpg|BK006934.2| 302036 - INS 
 tpg|BK006934.2| 52339 + tpg|BK006934.2| 51933 - INS 
 tpg|BK006934.2| 250454 + tpg|BK006934.2| 251156 - INS 
 tpg|BK006934.2| 82589 + tpg|BK006934.2| 81854 - INS 
 tpg|BK006934.2| 192879 + tpg|BK006934.2| 193363 - INS 
 tpg|BK006934.2| 16709 + tpg|BK006934.2| 16180 - INS 
 tpg|BK006934.2| 428931 + tpg|BK006934.2| 428451 - INS 
 tpg|BK006934.2| 26364 + tpg|BK006934.2| 26290 - INS 
 tpg|BK006934.2| 122910 + tpg|BK006934.2| 123051 - INS 
 tpg|BK006934.2| 77294 + tpg|BK006934.2| 77923 - INS 
 tpg|BK006934.2| 220134 + tpg|BK006934.2| 220611 - INS 
 tpg|BK006934.2| 365137 + tpg|BK006934.2| 365582 - INS 
 tpg|BK006934.2| 331780 + tpg|BK006934.2| 331522 - INS 
 tpg|BK006941.2| 770154 + tpg|BK006941.2| 769730 - INS 
 tpg|BK006934.2| 384066 + tpg|BK006934.2| 384465 - INS 
 tpg|BK006941.2| 627866 + tpg|BK006941.2| 627320 - INS 
 tpg|BK006934.2| 96634 + tpg|BK006934.2| 96460 - INS 
 tpg|BK006941.2| 55458 + tpg|BK006941.2| 54982 - INS 
 tpg|BK006934.2| 151116 + tpg|BK006934.2| 151326 - INS 
 tpg|BK006934.2| 520558 + tpg|BK006934.2| 520314 - INS 
 tpg|BK006934.2| 148358 + tpg|BK006934.2| 147883 - INS 
 tpg|BK006941.2| 379906 + tpg|BK006941.2| 379924 - INS 
 tpg|BK006934.2| 299748 + tpg|BK006934.2| 299320 - INS 
 tpg|BK006934.2| 273254 + tpg|BK006934.2| 273187 - INS 
 tpg|BK006934.2| 138558 + tpg|BK006934.2| 139330 - INS 
 tpg|BK006941.2| 654681 + tpg|BK006941.2| 655230 - INS 
 tpg|BK006934.2| 401277 + tpg|BK006934.2| 401062 - INS 
 tpg|BK006941.2| 197444 + tpg|BK006941.2| 197335 - INS 
 tpg|BK006934.2| 52884 + tpg|BK006934.2| 52917 - INS 
 tpg|BK006934.2| 242010 + tpg|BK006934.2| 241832 - INS 
 tpg|BK006934.2| 376430 + tpg|BK006934.2| 375973 - INS 
 tpg|BK006934.2| 38996 + tpg|BK006934.2| 38779 - INS 
 tpg|BK006941.2| 858959 + tpg|BK006941.2| 859122 - INS 
 tpg|BK006934.2| 219462 + tpg|BK006934.2| 219019 - INS 
 tpg|BK006934.2| 167345 + tpg|BK006934.2| 167013 - INS 
 tpg|BK006934.2| 199144 + tpg|BK006934.2| 198444 - INS 
 tpg|BK006941.2| 874739 + tpg|BK006941.2| 874873 - INS 
 tpg|BK006934.2| 493357 + tpg|BK006934.2| 493385 - INS 
 tpg|BK006934.2| 50898 + tpg|BK006934.2| 50981 - INS 
 tpg|BK006934.2| 310319 + tpg|BK006934.2| 310628 - INS 
 tpg|BK006941.2| 262219 + tpg|BK006941.2| 262110 - INS 
 tpg|BK006934.2| 434236 + tpg|BK006934.2| 434210 - INS 
 tpg|BK006934.2| 35127 + tpg|BK006934.2| 34970 - INS 
 tpg|BK006941.2| 893755 + tpg|BK006941.2| 893430 - INS 
 tpg|BK006934.2| 195406 + tpg|BK006934.2| 195023 - INS 
 tpg|BK006934.2| 53770 + tpg|BK006934.2| 54414 - INS 
 tpg|BK006934.2| 30152 + tpg|BK006934.2| 30559 - INS 
 tpg|BK006934.2| 359686 + tpg|BK006934.2| 359542 - INS 
 tpg|BK006941.2| 872950 + tpg|BK006941.2| 873644 - INS 
 tpg|BK006934.2| 414920 + tpg|BK006934.2| 414781 - INS 
 tpg|BK006934.2| 467960 + tpg|BK006934.2| 468178 - INS 
 tpg|BK006934.2| 212198 + tpg|BK006934.2| 212001 - INS 
 tpg|BK006934.2| 22113 + tpg|BK006934.2| 22028 - INS 
 tpg|BK006941.2| 484495 + tpg|BK006941.2| 484211 - INS 
 tpg|BK006934.2| 155869 + tpg|BK006934.2| 155268 - INS 
 tpg|BK006941.2| 304172 + tpg|BK006941.2| 303674 - INS 
 tpg|BK006934.2| 465119 + tpg|BK006934.2| 465027 - INS 
 tpg|BK006934.2| 311983 + tpg|BK006934.2| 311317 - INS 
 tpg|BK006934.2| 293467 + tpg|BK006934.2| 293036 - INS 
 tpg|BK006934.2| 291621 + tpg|BK006934.2| 291411 - INS 
 tpg|BK006934.2| 405546 + tpg|BK006934.2| 405039 - INS 
 tpg|BK006934.2| 146225 + tpg|BK006934.2| 145803 - INS 
 tpg|BK006934.2| 344721 + tpg|BK006934.2| 344791 - INS 
 tpg|BK006934.2| 46166 + tpg|BK006934.2| 46723 - INS 
 tpg|BK006941.2| 1065600 + tpg|BK006941.2| 1065059 - INS 
 tpg|BK006934.2| 347921 + tpg|BK006934.2| 347568 - INS 
 tpg|BK006934.2| 106114 + tpg|BK006934.2| 105939 - INS 
 tpg|BK006941.2| 247987 + tpg|BK006941.2| 248126 - INS 
 tpg|BK006934.2| 62842 + tpg|BK006934.2| 62493 - INS 
 tpg|BK006934.2| 149004 + tpg|BK006934.2| 149302 - INS 
 tpg|BK006934.2| 291978 + tpg|BK006934.2| 292400 - INS 
 tpg|BK006941.2| 747085 + tpg|BK006941.2| 747657 - INS 
 tpg|BK006934.2| 96087 + tpg|BK006934.2| 95318 - INS 
 tpg|BK006941.2| 270899 + tpg|BK006941.2| 271352 - INS 
 tpg|BK006934.2| 67280 + tpg|BK006934.2| 66755 - INS 
 tpg|BK006934.2| 257823 + tpg|BK006934.2| 257576 - INS 
 tpg|BK006934.2| 319739 + tpg|BK006934.2| 320124 - INS 
 tpg|BK006934.2| 358749 + tpg|BK006934.2| 358760 - INS 
 tpg|BK006941.2| 313936 + tpg|BK006941.2| 313172 - INS 
 tpg|BK006934.2| 108799 + tpg|BK006934.2| 109087 - INS 
 tpg|BK006934.2| 205558 + tpg|BK006934.2| 206083 - INS 
 tpg|BK006934.2| 380655 + tpg|BK006934.2| 380188 - INS 
 tpg|BK006941.2| 808815 + tpg|BK006941.2| 808403 - INS 
 tpg|BK006934.2| 353312 + tpg|BK006934.2| 353011 - INS 
 tpg|BK006941.2| 69083 + tpg|BK006941.2| 68827 - INS 
 tpg|BK006934.2| 356077 + tpg|BK006934.2| 355840 - INS 
 tpg|BK006934.2| 332722 + tpg|BK006934.2| 331959 - INS 
 tpg|BK006934.2| 503567 + tpg|BK006934.2| 504161 - INS 
 tpg|BK006941.2| 1583 + tpg|BK006941.2| 1085 - INS 
 tpg|BK006934.2| 425349 + tpg|BK006934.2| 424623 - INS 
 tpg|BK006934.2| 297634 + tpg|BK006934.2| 297572 - INS 
 tpg|BK006941.2| 640633 + tpg|BK006941.2| 640877 - INS 
 tpg|BK006934.2| 314936 + tpg|BK006934.2| 314871 - INS 
 tpg|BK006934.2| 339263 + tpg|BK006934.2| 339046 - INS 
 tpg|BK006934.2| 460796 + tpg|BK006934.2| 460035 - INS 
 tpg|BK006934.2| 370706 + tpg|BK006934.2| 370592 - INS 
 tpg|BK006934.2| 80043 + tpg|BK006934.2| 79983 - INS 
 tpg|BK006934.2| 525548 + tpg|BK006934.2| 524891 - INS 
 tpg|BK006941.2| 272982 + tpg|BK006941.2| 272573 - INS 
 tpg|BK006934.2| 294408 + tpg|BK006934.2| 293927 - INS 
 tpg|BK006934.2| 375831 + tpg|BK006934.2| 375134 - INS 
 tpg|BK006941.2| 267669 + tpg|BK006941.2| 267001 - INS 
 tpg|BK006934.2| 117153 + tpg|BK006934.2| 117450 - INS 
 tpg|BK006934.2| 137982 + tpg|BK006934.2| 137426 - INS 
 tpg|BK006934.2| 25433 + tpg|BK006934.2| 25614 - INS 
 tpg|BK006934.2| 473121 + tpg|BK006934.2| 473259 - INS 
 tpg|BK006934.2| 234678 + tpg|BK006934.2| 234714 - INS 
 tpg|BK006941.2| 242164 + tpg|BK006941.2| 241984 - INS 
 tpg|BK006934.2| 169627 + tpg|BK006934.2| 169679 - INS 
 tpg|BK006934.2| 103503 + tpg|BK006934.2| 102747 - INS 
 tpg|BK006934.2| 163780 + tpg|BK006934.2| 163719 - INS 
 tpg|BK006934.2| 24556 + tpg|BK006934.2| 24395 - INS 
 tpg|BK006934.2| 303595 + tpg|BK006934.2| 303302 - INS 
 tpg|BK006934.2| 150476 + tpg|BK006934.2| 150012 - INS 
 tpg|BK006941.2| 357662 + tpg|BK006941.2| 357625 - INS 
 tpg|BK006934.2| 278231 + tpg|BK006934.2| 278664 - INS 
 tpg|BK006941.2| 974777 + tpg|BK006941.2| 975549 - INS 
 tpg|BK006941.2| 420472 + tpg|BK006941.2| 420867 - INS 
 tpg|BK006934.2| 41185 + tpg|BK006934.2| 40623 - INS 
 tpg|BK006941.2| 733481 + tpg|BK006941.2| 733879 - INS 
 tpg|BK006934.2| 529603 + tpg|BK006934.2| 528873 - INS 
 tpg|BK006934.2| 521117 + tpg|BK006934.2| 520796 - INS 
 tpg|BK006941.2| 1061642 + tpg|BK006941.2| 1061796 - INS 
 tpg|BK006934.2| 485242 + tpg|BK006934.2| 485322 - INS 
 tpg|BK006934.2| 345769 + tpg|BK006934.2| 346231 - INS 
 tpg|BK006941.2| 511892 + tpg|BK006941.2| 511664 - INS 
 tpg|BK006934.2| 554635 + tpg|BK006934.2| 554962 - INS 
 tpg|BK006934.2| 202547 + tpg|BK006934.2| 202631 - INS 
 tpg|BK006934.2| 190406 + tpg|BK006934.2| 189962 - INS 
 tpg|BK006941.2| 833910 + tpg|BK006941.2| 833991 - INS 
 tpg|BK006934.2| 15095 + tpg|BK006934.2| 14969 - INS 
 tpg|BK006941.2| 979066 + tpg|BK006941.2| 978664 - INS 
 tpg|BK006934.2| 269140 + tpg|BK006934.2| 269546 - INS 
 tpg|BK006934.2| 455084 + tpg|BK006934.2| 454944 - INS 
 tpg|BK006934.2| 179078 + tpg|BK006934.2| 178956 - INS 
 tpg|BK006934.2| 431853 + tpg|BK006934.2| 431536 - INS 
 tpg|BK006934.2| 211084 + tpg|BK006934.2| 211262 - INS 
 tpg|BK006941.2| 447186 + tpg|BK006941.2| 447958 - INS 
 tpg|BK006934.2| 260934 + tpg|BK006934.2| 260376 - INS 
 tpg|BK006934.2| 510489 + tpg|BK006934.2| 510530 - INS GTG
 tpg|BK006941.2| 375847 + tpg|BK006941.2| 376156 - INS 
 tpg|BK006934.2| 492257 + tpg|BK006934.2| 492192 - INS 
 tpg|BK006934.2| 223088 + tpg|BK006934.2| 223307 - INS 
 tpg|BK006934.2| 229124 + tpg|BK006934.2| 229277 - INS 
 tpg|BK006934.2| 131971 + tpg|BK006934.2| 132495 - INS 
 tpg|BK006934.2| 531252 + tpg|BK006934.2| 530778 - INS 
 tpg|BK006941.2| 4615 + tpg|BK006941.2| 4679 - INS 
 tpg|BK006934.2| 448262 + tpg|BK006934.2| 448452 - INS 
 tpg|BK006934.2| 393341 + tpg|BK006934.2| 393386 - INS 
 tpg|BK006934.2| 398497 + tpg|BK006934.2| 398384 - INS 
 tpg|BK006941.2| 76720 + tpg|BK006941.2| 77127 - INS 
 tpg|BK006934.2| 233342 + tpg|BK006934.2| 232718 - INS 
 tpg|BK006934.2| 442615 + tpg|BK006934.2| 442550 - INS 
 tpg|BK006934.2| 425700 + tpg|BK006934.2| 425351 - INS 
 tpg|BK006934.2| 83305 + tpg|BK006934.2| 83213 - INS 
 tpg|BK006934.2| 303061 + tpg|BK006934.2| 302595 - INS 
 tpg|BK006934.2| 33039 + tpg|BK006934.2| 33132 - INS 
 tpg|BK006934.2| 305389 + tpg|BK006934.2| 305179 - INS 
 tpg|BK006934.2| 554081 + tpg|BK006934.2| 553393 - INS 
 tpg|BK006941.2| 732667 + tpg|BK006941.2| 733035 - INS 
 tpg|BK006941.2| 60469 + tpg|BK006941.2| 60952 - INS 
 tpg|BK006941.2| 851498 + tpg|BK006941.2| 851704 - INS 
 tpg|BK006934.2| 357631 + tpg|BK006934.2| 357219 - INS 
 tpg|BK006934.2| 156706 + tpg|BK006934.2| 156744 - INS 
 tpg|BK006934.2| 45148 + tpg|BK006934.2| 45495 - INS 
 tpg|BK006934.2| 187724 + tpg|BK006934.2| 187451 - INS 
 tpg|BK006941.2| 433936 + tpg|BK006941.2| 433883 - INS 
 tpg|BK006934.2| 309648 + tpg|BK006934.2| 309929 - INS 
 tpg|BK006934.2| 216987 + tpg|BK006934.2| 217241 - INS 
 tpg|BK006934.2| 527585 + tpg|BK006934.2| 527671 - INS 
 tpg|BK006934.2| 471201 + tpg|BK006934.2| 470963 - INS 
 tpg|BK006934.2| 254790 + tpg|BK006934.2| 254936 - INS 
 tpg|BK006934.2| 451748 + tpg|BK006934.2| 451321 - INS 
 tpg|BK006941.2| 102741 + tpg|BK006941.2| 102678 - INS ATATAGCTTAT
 tpg|BK006934.2| 27220 + tpg|BK006934.2| 27235 - INS 
 tpg|BK006934.2| 111464 + tpg|BK006934.2| 111121 - INS 
 tpg|BK006934.2| 373265 + tpg|BK006934.2| 372748 - INS 
 tpg|BK006934.2| 97059 + tpg|BK006934.2| 97676 - INS 
 tpg|BK006934.2| 521713 + tpg|BK006934.2| 521460 - INS 
 tpg|BK006934.2| 479829 + tpg|BK006934.2| 479666 - INS 
 tpg|BK006934.2| 427380 + tpg|BK006934.2| 426681 - INS 
 tpg|BK006934.2| 429373 + tpg|BK006934.2| 429263 - INS 
 tpg|BK006934.2| 336198 + tpg|BK006934.2| 335843 - INS 
 tpg|BK006934.2| 421532 + tpg|BK006934.2| 421421 - INS 
 tpg|BK006934.2| 108236 + tpg|BK006934.2| 108215 - INS 
 tpg|BK006934.2| 411071 + tpg|BK006934.2| 410784 - INS 
 tpg|BK006934.2| 388295 + tpg|BK006934.2| 388367 - INS 
 tpg|BK006934.2| 61636 + tpg|BK006934.2| 61387 - INS 
 tpg|BK006934.2| 28141 + tpg|BK006934.2| 27984 - INS 
 tpg|BK006934.2| 447573 + tpg|BK006934.2| 447925 - INS 
 tpg|BK006934.2| 336892 + tpg|BK006934.2| 336479 - INS 
 tpg|BK006934.2| 457325 + tpg|BK006934.2| 457266 - INS 
 tpg|BK006934.2| 85445 + tpg|BK006934.2| 85277 - INS 
 tpg|BK006934.2| 333067 + tpg|BK006934.2| 332876 - INS 
 tpg|BK006934.2| 348540 + tpg|BK006934.2| 348524 - INS 
 tpg|BK006941.2| 849219 + tpg|BK006941.2| 848540 - INS 
 tpg|BK006934.2| 476225 + tpg|BK006934.2| 476228 - INS 
 tpg|BK006934.2| 11968 + tpg|BK006934.2| 12224 - INS 
 tpg|BK006934.2| 287507 + tpg|BK006934.2| 287008 - INS 
 tpg|BK006941.2| 236258 + tpg|BK006941.2| 236484 - INS 
 tpg|BK006934.2| 67753 + tpg|BK006934.2| 68069 - INS 
 tpg|BK006934.2| 206988 + tpg|BK006934.2| 207225 - INS 
 tpg|BK006934.2| 494766 + tpg|BK006934.2| 494549 - INS 
 tpg|BK006934.2| 502838 + tpg|BK006934.2| 502741 - INS 
 tpg|BK006941.2| 363239 + tpg|BK006941.2| 362820 - INS 
 tpg|BK006941.2| 930563 + tpg|BK006941.2| 930075 - INS 
 tpg|BK006934.2| 167916 + tpg|BK006934.2| 168057 - INS 
 tpg|BK006934.2| 274221 + tpg|BK006934.2| 273681 - INS 
 tpg|BK006934.2| 72425 + tpg|BK006934.2| 72469 - INS 
 tpg|BK006934.2| 270644 + tpg|BK006934.2| 270298 - INS 
 tpg|BK006941.2| 372866 + tpg|BK006941.2| 372743 - INS 
 tpg|BK006934.2| 484538 + tpg|BK006934.2| 484225 - INS 
 tpg|BK006934.2| 260122 + tpg|BK006934.2| 259690 - INS 
 tpg|BK006934.2| 349723 + tpg|BK006934.2| 349582 - INS 
 tpg|BK006934.2| 340752 + tpg|BK006934.2| 340976 - INS 
 tpg|BK006941.2| 510610 + tpg|BK006941.2| 510319 - INS 
 tpg|BK006934.2| 258581 + tpg|BK006934.2| 259109 - INS 
 tpg|BK006934.2| 300218 + tpg|BK006934.2| 300654 - INS 
 tpg|BK006934.2| 524983 + tpg|BK006934.2| 524432 - INS 
 tpg|BK006934.2| 172089 + tpg|BK006934.2| 172025 - INS 
 tpg|BK006934.2| 65724 + tpg|BK006934.2| 65426 - INS 
 tpg|BK006934.2| 329012 + tpg|BK006934.2| 329490 - INS 
 tpg|BK006934.2| 233589 + tpg|BK006934.2| 234211 - INS 
 tpg|BK006941.2| 892441 + tpg|BK006941.2| 892585 - INS 
 tpg|BK006941.2| 79348 + tpg|BK006941.2| 79746 - INS 
 tpg|BK006941.2| 96506 + tpg|BK006941.2| 95999 - INS 
 tpg|BK006941.2| 805085 + tpg|BK006941.2| 804586 - INS 
 tpg|BK006941.2| 126367 + tpg|BK006941.2| 126279 - INS 
 tpg|BK006941.2| 140315 + tpg|BK006941.2| 140338 - INS 
 tpg|BK006941.2| 411084 + tpg|BK006941.2| 410780 - INS 
 tpg|BK006941.2| 850034 + tpg|BK006941.2| 849510 - INS 
 tpg|BK006941.2| 993425 + tpg|BK006941.2| 992791 - INS 
 tpg|BK006941.2| 414804 + tpg|BK006941.2| 414054 - INS 
 tpg|BK006941.2| 899035 + tpg|BK006941.2| 898660 - INS 
 tpg|BK006941.2| 352175 + tpg|BK006941.2| 351752 - INS 
 tpg|BK006941.2| 397794 + tpg|BK006941.2| 398044 - INS 
 tpg|BK006941.2| 268687 + tpg|BK006941.2| 268832 - INS 
 tpg|BK006941.2| 593274 + tpg|BK006941.2| 593037 - INS 
 tpg|BK006941.2| 643324 + tpg|BK006941.2| 643168 - INS 
 tpg|BK006941.2| 625919 + tpg|BK006941.2| 625731 - INS 
 tpg|BK006941.2| 666849 + tpg|BK006941.2| 667499 - INS 
 tpg|BK006941.2| 58553 + tpg|BK006941.2| 57922 - INS 
 tpg|BK006941.2| 224643 + tpg|BK006941.2| 224929 - INS 
 tpg|BK006941.2| 134594 + tpg|BK006941.2| 134843 - INS 
 tpg|BK006941.2| 352758 + tpg|BK006941.2| 352989 - INS 
 tpg|BK006941.2| 783752 + tpg|BK006941.2| 783382 - INS 
 tpg|BK006941.2| 885858 + tpg|BK006941.2| 885856 - INS 
 tpg|BK006941.2| 927408 + tpg|BK006941.2| 927125 - INS 
 tpg|BK006941.2| 476034 + tpg|BK006941.2| 476594 - INS 
 tpg|BK006941.2| 943143 + tpg|BK006941.2| 942701 - INS 
 tpg|BK006941.2| 501846 + tpg|BK006941.2| 501413 - INS 
 tpg|BK006941.2| 679070 + tpg|BK006941.2| 678876 - INS 
 tpg|BK006941.2| 547453 + tpg|BK006941.2| 547243 - INS 
 tpg|BK006941.2| 624392 + tpg|BK006941.2| 623723 - INS 
 tpg|BK006941.2| 1071244 + tpg|BK006941.2| 1070769 - INS 
 tpg|BK006941.2| 405607 + tpg|BK006941.2| 406160 - INS 
 tpg|BK006941.2| 828869 + tpg|BK006941.2| 828254 - INS 
 tpg|BK006941.2| 196506 + tpg|BK006941.2| 195810 - INS 
 tpg|BK006941.2| 199311 + tpg|BK006941.2| 199164 - INS 
 tpg|BK006941.2| 448387 + tpg|BK006941.2| 448560 - INS 
 tpg|BK006941.2| 956394 + tpg|BK006941.2| 956040 - INS 
 tpg|BK006941.2| 1049329 + tpg|BK006941.2| 1049416 - INS 
 tpg|BK006941.2| 350400 + tpg|BK006941.2| 349718 - INS 
 tpg|BK006941.2| 991885 + tpg|BK006941.2| 991112 - INS 
 tpg|BK006941.2| 1012280 + tpg|BK006941.2| 1011881 - INS TAACCATGAGACAA
 tpg|BK006941.2| 188338 + tpg|BK006941.2| 188047 - INS 
 tpg|BK006941.2| 577132 + tpg|BK006941.2| 576621 - INS 
 tpg|BK006941.2| 297499 + tpg|BK006941.2| 297958 - INS 
 tpg|BK006941.2| 453899 + tpg|BK006941.2| 453333 - INS 
 tpg|BK006941.2| 911405 + tpg|BK006941.2| 910909 - INS 
 tpg|BK006941.2| 124228 + tpg|BK006941.2| 124044 - INS 
 tpg|BK006941.2| 598326 + tpg|BK006941.2| 597791 - INS 
 tpg|BK006941.2| 578044 + tpg|BK006941.2| 578742 - INS 
 tpg|BK006941.2| 74400 + tpg|BK006941.2| 74400 - INS 
 tpg|BK006941.2| 440845 + tpg|BK006941.2| 440383 - INS 
 tpg|BK006941.2| 5485 + tpg|BK006941.2| 5517 - INS 
 tpg|BK006941.2| 261002 + tpg|BK006941.2| 260372 - INS 
 tpg|BK006941.2| 672817 + tpg|BK006941.2| 672255 - INS 
 tpg|BK006941.2| 192810 + tpg|BK006941.2| 192051 - INS 
 tpg|BK006941.2| 384366 + tpg|BK006941.2| 384238 - INS 
 tpg|BK006941.2| 204380 + tpg|BK006941.2| 203799 - INS 
 tpg|BK006941.2| 443286 + tpg|BK006941.2| 443270 - INS 
 tpg|BK006941.2| 426928 + tpg|BK006941.2| 426778 - INS 
 tpg|BK006941.2| 116700 + tpg|BK006941.2| 115963 - INS 
 tpg|BK006941.2| 81054 + tpg|BK006941.2| 81316 - INS 
 tpg|BK006941.2| 233039 + tpg|BK006941.2| 232468 - INS 
 tpg|BK006941.2| 395706 + tpg|BK006941.2| 395199 - INS 
 tpg|BK006941.2| 857057 + tpg|BK006941.2| 856965 - INS 
 tpg|BK006938.2| 1247245 + tpg|BK006938.2| 1247135 - INS 
 tpg|BK006941.2| 968228 + tpg|BK006941.2| 967744 - INS 
 tpg|BK006938.2| 147581 + tpg|BK006938.2| 147605 - INS 
 tpg|BK006941.2| 39726 + tpg|BK006941.2| 39722 - INS 
 tpg|BK006941.2| 504314 + tpg|BK006941.2| 503781 - INS 
 tpg|BK006941.2| 341895 + tpg|BK006941.2| 342414 - INS 
 tpg|BK006938.2| 451323 + tpg|BK006938.2| 450887 - INS 
 tpg|BK006941.2| 187664 + tpg|BK006941.2| 187320 - INS 
 tpg|BK006941.2| 339412 + tpg|BK006941.2| 339164 - INS 
 tpg|BK006938.2| 384811 + tpg|BK006938.2| 385099 - INS 
 tpg|BK006941.2| 1053019 + tpg|BK006941.2| 1052823 - INS 
 tpg|BK006941.2| 321505 + tpg|BK006941.2| 321559 - INS 
 tpg|BK006941.2| 636152 + tpg|BK006941.2| 636564 - INS 
 tpg|BK006941.2| 301891 + tpg|BK006941.2| 301721 - INS 
 tpg|BK006941.2| 291382 + tpg|BK006941.2| 290802 - INS 
 tpg|BK006938.2| 411659 + tpg|BK006938.2| 411552 - INS 
 tpg|BK006938.2| 1227144 + tpg|BK006938.2| 1226873 - INS 
 tpg|BK006941.2| 534167 + tpg|BK006941.2| 534471 - INS 
 tpg|BK006938.2| 1431911 + tpg|BK006938.2| 1432307 - INS 
 tpg|BK006941.2| 181500 + tpg|BK006941.2| 180995 - INS 
 tpg|BK006941.2| 845065 + tpg|BK006941.2| 845170 - INS 
 tpg|BK006941.2| 148885 + tpg|BK006941.2| 149093 - INS 
 tpg|BK006941.2| 26652 + tpg|BK006941.2| 26942 - INS 
 tpg|BK006938.2| 406301 + tpg|BK006938.2| 407040 - INS 
 tpg|BK006941.2| 998377 + tpg|BK006941.2| 998432 - INS 
 tpg|BK006941.2| 10182 + tpg|BK006941.2| 9786 - INS 
 tpg|BK006938.2| 105424 + tpg|BK006938.2| 105752 - INS 
 tpg|BK006941.2| 390001 + tpg|BK006941.2| 389728 - INS 
 tpg|BK006941.2| 915426 + tpg|BK006941.2| 915566 - INS 
 tpg|BK006941.2| 380344 + tpg|BK006941.2| 381022 - INS 
 tpg|BK006941.2| 97757 + tpg|BK006941.2| 98163 - INS 
 tpg|BK006941.2| 824017 + tpg|BK006941.2| 823446 - INS 
 tpg|BK006941.2| 360180 + tpg|BK006941.2| 360321 - INS 
 tpg|BK006941.2| 866722 + tpg|BK006941.2| 866680 - INS 
 tpg|BK006938.2| 1525161 + tpg|BK006938.2| 1524611 - INS 
 tpg|BK006941.2| 156905 + tpg|BK006941.2| 156984 - INS 
 tpg|BK006938.2| 1059242 + tpg|BK006938.2| 1058899 - INS 
 tpg|BK006941.2| 454619 + tpg|BK006941.2| 453974 - INS 
 tpg|BK006941.2| 741567 + tpg|BK006941.2| 741045 - INS 
 tpg|BK006941.2| 200255 + tpg|BK006941.2| 200573 - INS 
 tpg|BK006941.2| 551357 + tpg|BK006941.2| 550684 - INS 
 tpg|BK006941.2| 170959 + tpg|BK006941.2| 170657 - INS 
 tpg|BK006941.2| 1053881 + tpg|BK006941.2| 1053498 - INS 
 tpg|BK006941.2| 1044943 + tpg|BK006941.2| 1044714 - INS 
 tpg|BK006941.2| 976698 + tpg|BK006941.2| 977336 - INS 
 tpg|BK006941.2| 1005367 + tpg|BK006941.2| 1005356 - INS 
 tpg|BK006941.2| 190787 + tpg|BK006941.2| 190125 - INS 
 tpg|BK006941.2| 520659 + tpg|BK006941.2| 521104 - INS 
 tpg|BK006941.2| 198473 + tpg|BK006941.2| 198299 - INS 
 tpg|BK006941.2| 962757 + tpg|BK006941.2| 962358 - INS 
 tpg|BK006941.2| 762233 + tpg|BK006941.2| 762393 - INS 
 tpg|BK006941.2| 1057257 + tpg|BK006941.2| 1057253 - INS 
 tpg|BK006941.2| 418161 + tpg|BK006941.2| 418119 - INS 
 tpg|BK006941.2| 799737 + tpg|BK006941.2| 799783 - INS 
 tpg|BK006941.2| 588124 + tpg|BK006941.2| 587642 - INS 
 tpg|BK006941.2| 336194 + tpg|BK006941.2| 336526 - INS 
 tpg|BK006941.2| 864691 + tpg|BK006941.2| 864728 - INS 
 tpg|BK006941.2| 1050869 + tpg|BK006941.2| 1051261 - INS 
 tpg|BK006941.2| 948910 + tpg|BK006941.2| 948851 - INS 
 tpg|BK006941.2| 292178 + tpg|BK006941.2| 292318 - INS 
 tpg|BK006941.2| 757813 + tpg|BK006941.2| 757141 - INS 
 tpg|BK006941.2| 786060 + tpg|BK006941.2| 785700 - INS 
 tpg|BK006941.2| 78513 + tpg|BK006941.2| 78391 - INS 
 tpg|BK006941.2| 371225 + tpg|BK006941.2| 370957 - INS 
 tpg|BK006941.2| 950108 + tpg|BK006941.2| 950034 - INS 
 tpg|BK006941.2| 963562 + tpg|BK006941.2| 963466 - INS 
 tpg|BK006941.2| 343416 + tpg|BK006941.2| 344143 - INS 
 tpg|BK006941.2| 980682 + tpg|BK006941.2| 979934 - INS 
 tpg|BK006941.2| 305744 + tpg|BK006941.2| 305188 - INS 
 tpg|BK006941.2| 1047543 + tpg|BK006941.2| 1047145 - INS 
 tpg|BK006941.2| 590842 + tpg|BK006941.2| 591262 - INS 
 tpg|BK006941.2| 602952 + tpg|BK006941.2| 602224 - INS 
 tpg|BK006941.2| 184813 + tpg|BK006941.2| 184684 - INS 
 tpg|BK006941.2| 925157 + tpg|BK006941.2| 924514 - INS 
 tpg|BK006941.2| 856110 + tpg|BK006941.2| 855570 - INS 
 tpg|BK006941.2| 790491 + tpg|BK006941.2| 789940 - INS 
 tpg|BK006941.2| 76045 + tpg|BK006941.2| 75809 - INS 
 tpg|BK006941.2| 104810 + tpg|BK006941.2| 104583 - INS 
 tpg|BK006941.2| 211364 + tpg|BK006941.2| 211673 - INS 
 tpg|BK006941.2| 746209 + tpg|BK006941.2| 745977 - INS 
 tpg|BK006941.2| 378771 + tpg|BK006941.2| 378080 - INS 
 tpg|BK006941.2| 941648 + tpg|BK006941.2| 941603 - INS 
 tpg|BK006941.2| 697928 + tpg|BK006941.2| 697505 - INS 
 tpg|BK006938.2| 91496 + tpg|BK006938.2| 92270 - INS 
 tpg|BK006941.2| 127756 + tpg|BK006941.2| 128375 - INS 
 tpg|BK006941.2| 676435 + tpg|BK006941.2| 676472 - INS 
 tpg|BK006938.2| 408776 + tpg|BK006938.2| 408882 - INS 
 tpg|BK006941.2| 983676 + tpg|BK006941.2| 983403 - INS 
 tpg|BK006941.2| 527405 + tpg|BK006941.2| 526815 - INS 
 tpg|BK006941.2| 328186 + tpg|BK006941.2| 327739 - INS 
 tpg|BK006941.2| 24426 + tpg|BK006941.2| 23969 - INS 
 tpg|BK006941.2| 599997 + tpg|BK006941.2| 600161 - INS 
 tpg|BK006941.2| 1010649 + tpg|BK006941.2| 1010052 - INS 
 tpg|BK006938.2| 652804 + tpg|BK006938.2| 652634 - INS 
 tpg|BK006941.2| 273787 + tpg|BK006941.2| 273223 - INS 
 tpg|BK006938.2| 67621 + tpg|BK006938.2| 67147 - INS 
 tpg|BK006941.2| 1013682 + tpg|BK006941.2| 1013301 - INS 
 tpg|BK006941.2| 287101 + tpg|BK006941.2| 286676 - INS 
 tpg|BK006941.2| 672422 + tpg|BK006941.2| 671756 - INS 
 tpg|BK006938.2| 485177 + tpg|BK006938.2| 485572 - INS 
 tpg|BK006938.2| 677805 + tpg|BK006938.2| 678093 - INS 
 tpg|BK006938.2| 1078043 + tpg|BK006938.2| 1078098 - INS 
 tpg|BK006941.2| 586616 + tpg|BK006941.2| 586999 - INS 
 tpg|BK006941.2| 492942 + tpg|BK006941.2| 492625 - INS 
 tpg|BK006941.2| 996095 + tpg|BK006941.2| 995479 - INS 
 tpg|BK006941.2| 43082 + tpg|BK006941.2| 42335 - INS 
 tpg|BK006938.2| 487458 + tpg|BK006938.2| 487331 - INS 
 tpg|BK006941.2| 461899 + tpg|BK006941.2| 461412 - INS 
 tpg|BK006941.2| 869929 + tpg|BK006941.2| 870046 - INS 
 tpg|BK006941.2| 879056 + tpg|BK006941.2| 878805 - INS 
 tpg|BK006941.2| 879631 + tpg|BK006941.2| 880317 - INS 
 tpg|BK006938.2| 573125 + tpg|BK006938.2| 572517 - INS 
 tpg|BK006938.2| 829106 + tpg|BK006938.2| 829317 - INS 
 tpg|BK006941.2| 260152 + tpg|BK006941.2| 259652 - INS 
 tpg|BK006938.2| 1341643 + tpg|BK006938.2| 1340913 - INS 
 tpg|BK006941.2| 147427 + tpg|BK006941.2| 147199 - INS 
 tpg|BK006938.2| 1188159 + tpg|BK006938.2| 1188685 - INS 
 tpg|BK006941.2| 641781 + tpg|BK006941.2| 641840 - INS 
 tpg|BK006941.2| 1041105 + tpg|BK006941.2| 1040331 - INS 
 tpg|BK006941.2| 499448 + tpg|BK006941.2| 499474 - INS 
 tpg|BK006941.2| 348660 + tpg|BK006941.2| 348290 - INS 
 tpg|BK006938.2| 464576 + tpg|BK006938.2| 463983 - INS 
 tpg|BK006941.2| 1069558 + tpg|BK006941.2| 1069243 - INS 
 tpg|BK006941.2| 763590 + tpg|BK006941.2| 763161 - INS 
 tpg|BK006938.2| 802363 + tpg|BK006938.2| 801604 - INS 
 tpg|BK006941.2| 796535 + tpg|BK006941.2| 796388 - INS 
 tpg|BK006941.2| 652765 + tpg|BK006941.2| 652551 - INS 
 tpg|BK006941.2| 127306 + tpg|BK006941.2| 127040 - INS 
 tpg|BK006941.2| 1079021 + tpg|BK006941.2| 1078312 - INS 
 tpg|BK006938.2| 108726 + tpg|BK006938.2| 108680 - INS 
 tpg|BK006938.2| 658565 + tpg|BK006938.2| 658178 - INS 
 tpg|BK006941.2| 54787 + tpg|BK006941.2| 54157 - INS 
 tpg|BK006941.2| 307981 + tpg|BK006941.2| 307426 - INS 
 tpg|BK006938.2| 859204 + tpg|BK006938.2| 859241 - INS 
 tpg|BK006941.2| 939424 + tpg|BK006941.2| 938963 - INS 
 tpg|BK006938.2| 699124 + tpg|BK006938.2| 698720 - INS 
 tpg|BK006941.2| 777470 + tpg|BK006941.2| 777599 - INS 
 tpg|BK006941.2| 677300 + tpg|BK006941.2| 677267 - INS 
 tpg|BK006941.2| 678099 + tpg|BK006941.2| 678554 - INS 
 tpg|BK006938.2| 1146120 + tpg|BK006938.2| 1145873 - INS 
 tpg|BK006941.2| 451959 + tpg|BK006941.2| 452411 - INS 
 tpg|BK006938.2| 975041 + tpg|BK006938.2| 974453 - INS 
 tpg|BK006941.2| 723041 + tpg|BK006941.2| 723262 - INS 
 tpg|BK006941.2| 398999 + tpg|BK006941.2| 398545 - INS 
 tpg|BK006938.2| 770153 + tpg|BK006938.2| 770627 - INS 
 tpg|BK006941.2| 402632 + tpg|BK006941.2| 402502 - INS 
 tpg|BK006938.2| 360187 + tpg|BK006938.2| 359761 - INS 
 tpg|BK006941.2| 115139 + tpg|BK006941.2| 114939 - INS 
 tpg|BK006941.2| 445150 + tpg|BK006941.2| 445449 - INS 
 tpg|BK006938.2| 258739 + tpg|BK006938.2| 258846 - INS 
 tpg|BK006941.2| 761316 + tpg|BK006941.2| 761674 - INS 
 tpg|BK006938.2| 272280 + tpg|BK006938.2| 272547 - INS 
 tpg|BK006941.2| 839441 + tpg|BK006941.2| 839260 - INS 
 tpg|BK006941.2| 840167 + tpg|BK006941.2| 839885 - INS 
 tpg|BK006941.2| 408312 + tpg|BK006941.2| 407833 - INS 
 tpg|BK006938.2| 686442 + tpg|BK006938.2| 685845 - INS 
 tpg|BK006941.2| 841224 + tpg|BK006941.2| 841316 - INS 
 tpg|BK006941.2| 63937 + tpg|BK006941.2| 63521 - INS 
 tpg|BK006938.2| 1085456 + tpg|BK006938.2| 1085440 - INS 
 tpg|BK006941.2| 258019 + tpg|BK006941.2| 258754 - INS 
 tpg|BK006938.2| 113372 + tpg|BK006938.2| 113283 - INS 
 tpg|BK006941.2| 1001493 + tpg|BK006941.2| 1002265 - INS 
 tpg|BK006941.2| 13090 + tpg|BK006941.2| 13056 - INS 
 tpg|BK006938.2| 199059 + tpg|BK006938.2| 198923 - INS 
 tpg|BK006941.2| 524768 + tpg|BK006941.2| 524193 - INS 
 tpg|BK006941.2| 283256 + tpg|BK006941.2| 282704 - INS 
 tpg|BK006941.2| 1084285 + tpg|BK006941.2| 1083981 - INS 
 tpg|BK006941.2| 358693 + tpg|BK006941.2| 359297 - INS 
 tpg|BK006941.2| 1060584 + tpg|BK006941.2| 1060033 - INS 
 tpg|BK006941.2| 1058288 + tpg|BK006941.2| 1058242 - INS 
 tpg|BK006941.2| 548049 + tpg|BK006941.2| 548183 - INS 
 tpg|BK006938.2| 1521151 + tpg|BK006938.2| 1521756 - INS 
 tpg|BK006938.2| 1081967 + tpg|BK006938.2| 1081772 - INS 
 tpg|BK006941.2| 1034665 + tpg|BK006941.2| 1034142 - INS 
 tpg|BK006941.2| 264957 + tpg|BK006941.2| 264672 - INS 
 tpg|BK006938.2| 868652 + tpg|BK006938.2| 868183 - INS 
 tpg|BK006941.2| 304943 + tpg|BK006941.2| 304669 - INS 
 tpg|BK006938.2| 605344 + tpg|BK006938.2| 604600 - INS 
 tpg|BK006941.2| 186020 + tpg|BK006941.2| 185586 - INS 
 tpg|BK006941.2| 165369 + tpg|BK006941.2| 166124 - INS 
 tpg|BK006938.2| 703215 + tpg|BK006938.2| 702618 - INS 
 tpg|BK006941.2| 584546 + tpg|BK006941.2| 583777 - INS 
 tpg|BK006938.2| 954459 + tpg|BK006938.2| 954222 - INS 
 tpg|BK006941.2| 732005 + tpg|BK006941.2| 731826 - INS 
 tpg|BK006938.2| 141182 + tpg|BK006938.2| 141786 - INS 
 tpg|BK006941.2| 620710 + tpg|BK006941.2| 620146 - INS 
 tpg|BK006938.2| 1281991 + tpg|BK006938.2| 1282523 - INS 
 tpg|BK006941.2| 734945 + tpg|BK006941.2| 734731 - INS 
 tpg|BK006941.2| 971681 + tpg|BK006941.2| 971338 - INS 
 tpg|BK006938.2| 1344628 + tpg|BK006938.2| 1343997 - INS 
 tpg|BK006941.2| 144239 + tpg|BK006941.2| 144509 - INS 
 tpg|BK006938.2| 585234 + tpg|BK006938.2| 584758 - INS 
 tpg|BK006941.2| 543112 + tpg|BK006941.2| 543331 - INS 
 tpg|BK006941.2| 138392 + tpg|BK006941.2| 137834 - INS 
 tpg|BK006938.2| 146789 + tpg|BK006938.2| 147139 - INS 
 tpg|BK006941.2| 215030 + tpg|BK006941.2| 214883 - INS 
 tpg|BK006938.2| 282697 + tpg|BK006938.2| 282524 - INS 
 tpg|BK006938.2| 850242 + tpg|BK006938.2| 850790 - INS 
 tpg|BK006940.2| 159901 + tpg|BK006940.2| 159502 - INS 
 tpg|BK006938.2| 568122 + tpg|BK006938.2| 568200 - INS 
 tpg|BK006938.2| 297001 + tpg|BK006938.2| 296790 - INS 
 tpg|BK006938.2| 1441090 + tpg|BK006938.2| 1440789 - INS 
 tpg|BK006940.2| 65907 + tpg|BK006940.2| 65274 - INS 
 tpg|BK006941.2| 101480 + tpg|BK006941.2| 101274 - INS 
 tpg|BK006938.2| 319620 + tpg|BK006938.2| 319259 - INS 
 tpg|BK006941.2| 910104 + tpg|BK006941.2| 910169 - INS 
 tpg|BK006940.2| 123133 + tpg|BK006940.2| 123185 - INS 
 tpg|BK006941.2| 860749 + tpg|BK006941.2| 860102 - INS 
 tpg|BK006938.2| 39739 + tpg|BK006938.2| 39920 - INS 
 tpg|BK006941.2| 401418 + tpg|BK006941.2| 400963 - INS 
 tpg|BK006940.2| 182682 + tpg|BK006940.2| 182268 - INS 
 tpg|BK006941.2| 759624 + tpg|BK006941.2| 759592 - INS 
 tpg|BK006938.2| 1075444 + tpg|BK006938.2| 1075096 - INS 
 tpg|BK006941.2| 616800 + tpg|BK006941.2| 616254 - INS 
 tpg|BK006938.2| 555177 + tpg|BK006938.2| 554768 - INS 
 tpg|BK006940.2| 224612 + tpg|BK006940.2| 224592 - INS 
 tpg|BK006938.2| 246714 + tpg|BK006938.2| 246430 - INS 
 tpg|BK006940.2| 79852 + tpg|BK006940.2| 80255 - INS 
 tpg|BK006938.2| 525207 + tpg|BK006938.2| 524501 - INS 
 tpg|BK006941.2| 162935 + tpg|BK006941.2| 162450 - INS 
 tpg|BK006941.2| 438846 + tpg|BK006941.2| 439171 - INS 
 tpg|BK006940.2| 49557 + tpg|BK006940.2| 49719 - INS 
 tpg|BK006941.2| 656166 + tpg|BK006941.2| 656005 - INS 
 tpg|BK006938.2| 1193635 + tpg|BK006938.2| 1193466 - INS 
 tpg|BK006941.2| 546213 + tpg|BK006941.2| 545856 - INS 
 tpg|BK006940.2| 181161 + tpg|BK006940.2| 181267 - INS 
 tpg|BK006941.2| 997115 + tpg|BK006941.2| 997714 - INS 
 tpg|BK006938.2| 218992 + tpg|BK006938.2| 218504 - INS 
 tpg|BK006941.2| 1000326 + tpg|BK006941.2| 999963 - INS 
 tpg|BK006938.2| 1279438 + tpg|BK006938.2| 1278839 - INS 
 tpg|BK006941.2| 613902 + tpg|BK006941.2| 614217 - INS 
 tpg|BK006938.2| 53704 + tpg|BK006938.2| 53615 - INS 
 tpg|BK006940.2| 225920 + tpg|BK006940.2| 225571 - INS 
 tpg|BK006941.2| 586006 + tpg|BK006941.2| 585323 - INS 
 tpg|BK006938.2| 614070 + tpg|BK006938.2| 613690 - INS 
 tpg|BK006940.2| 205949 + tpg|BK006940.2| 205773 - INS 
 tpg|BK006941.2| 412549 + tpg|BK006941.2| 412178 - INS 
 tpg|BK006938.2| 906522 + tpg|BK006938.2| 906518 - INS 
 tpg|BK006941.2| 112556 + tpg|BK006941.2| 112755 - INS 
 tpg|BK006940.2| 90041 + tpg|BK006940.2| 90138 - INS 
 tpg|BK006938.2| 842323 + tpg|BK006938.2| 841633 - INS 
 tpg|BK006940.2| 87933 + tpg|BK006940.2| 87593 - INS 
 tpg|BK006938.2| 1261680 + tpg|BK006938.2| 1261130 - INS 
 tpg|BK006940.2| 254282 + tpg|BK006940.2| 254177 - INS 
 tpg|BK006940.2| 91625 + tpg|BK006940.2| 92322 - INS 
 tpg|BK006938.2| 229356 + tpg|BK006938.2| 229174 - INS 
 tpg|BK006940.2| 100952 + tpg|BK006940.2| 100451 - INS 
 tpg|BK006940.2| 110729 + tpg|BK006940.2| 111168 - INS 
 tpg|BK006941.2| 229552 + tpg|BK006941.2| 230135 - INS 
 tpg|BK006938.2| 150319 + tpg|BK006938.2| 150192 - INS 
 tpg|BK006940.2| 23768 + tpg|BK006940.2| 24095 - INS 
 tpg|BK006940.2| 168900 + tpg|BK006940.2| 168243 - INS 
 tpg|BK006941.2| 901339 + tpg|BK006941.2| 901434 - INS 
 tpg|BK006940.2| 154493 + tpg|BK006940.2| 154950 - INS 
 tpg|BK006941.2| 49934 + tpg|BK006941.2| 49211 - INS 
 tpg|BK006941.2| 430474 + tpg|BK006941.2| 430332 - INS 
 tpg|BK006940.2| 5538 + tpg|BK006940.2| 5465 - INS 
 tpg|BK006941.2| 84894 + tpg|BK006941.2| 84692 - INS 
 tpg|BK006941.2| 424204 + tpg|BK006941.2| 424199 - INS 
 tpg|BK006938.2| 86572 + tpg|BK006938.2| 86353 - INS 
 tpg|BK006940.2| 190153 + tpg|BK006940.2| 189725 - INS 
 tpg|BK006941.2| 82509 + tpg|BK006941.2| 82141 - INS 
 tpg|BK006940.2| 217226 + tpg|BK006940.2| 217611 - INS 
 tpg|BK006938.2| 413945 + tpg|BK006938.2| 413728 - INS 
 tpg|BK006941.2| 73297 + tpg|BK006941.2| 72692 - INS 
 tpg|BK006938.2| 1296077 + tpg|BK006938.2| 1296361 - INS 
 tpg|BK006940.2| 58607 + tpg|BK006940.2| 58397 - INS 
 tpg|BK006940.2| 165211 + tpg|BK006940.2| 164900 - INS 
 tpg|BK006941.2| 559119 + tpg|BK006941.2| 559078 - INS 
 tpg|BK006938.2| 1016886 + tpg|BK006938.2| 1016555 - INS 
 tpg|BK006940.2| 211415 + tpg|BK006940.2| 210861 - INS 
 tpg|BK006941.2| 743029 + tpg|BK006941.2| 743440 - INS 
 tpg|BK006938.2| 1003102 + tpg|BK006938.2| 1003835 - INS 
 tpg|BK006940.2| 93952 + tpg|BK006940.2| 94051 - INS 
 tpg|BK006941.2| 279590 + tpg|BK006941.2| 279054 - INS 
 tpg|BK006941.2| 284200 + tpg|BK006941.2| 284827 - INS 
 tpg|BK006940.2| 242305 + tpg|BK006940.2| 242303 - INS 
 tpg|BK006938.2| 1387237 + tpg|BK006938.2| 1387956 - INS 
 tpg|BK006941.2| 28054 + tpg|BK006941.2| 28623 - INS 
 tpg|BK006941.2| 9425 + tpg|BK006941.2| 8903 - INS 
 tpg|BK006941.2| 621942 + tpg|BK006941.2| 622330 - INS 
 tpg|BK006938.2| 560059 + tpg|BK006938.2| 560404 - INS 
 tpg|BK006940.2| 128240 + tpg|BK006940.2| 127735 - INS 
 tpg|BK006941.2| 1030664 + tpg|BK006941.2| 1031135 - INS 
 tpg|BK006940.2| 119390 + tpg|BK006940.2| 119427 - INS 
 tpg|BK006940.2| 246707 + tpg|BK006940.2| 246707 - INS 
 tpg|BK006938.2| 725324 + tpg|BK006938.2| 725717 - INS 
 tpg|BK006941.2| 515503 + tpg|BK006941.2| 515217 - INS ACGA
 tpg|BK006938.2| 18435 + tpg|BK006938.2| 18988 - INS 
 tpg|BK006940.2| 116999 + tpg|BK006940.2| 117021 - INS 
 tpg|BK006938.2| 126558 + tpg|BK006938.2| 126805 - INS 
 tpg|BK006941.2| 670045 + tpg|BK006941.2| 669633 - INS 
 tpg|BK006941.2| 133885 + tpg|BK006941.2| 133459 - INS 
 tpg|BK006940.2| 183420 + tpg|BK006940.2| 183650 - INS 
 tpg|BK006938.2| 131912 + tpg|BK006938.2| 131146 - INS 
 tpg|BK006941.2| 507650 + tpg|BK006941.2| 507167 - INS 
 tpg|BK006941.2| 730154 + tpg|BK006941.2| 730411 - INS 
 tpg|BK006938.2| 1318393 + tpg|BK006938.2| 1318627 - INS 
 tpg|BK006941.2| 346708 + tpg|BK006941.2| 346533 - INS 
 tpg|BK006938.2| 1383220 + tpg|BK006938.2| 1382550 - INS 
 tpg|BK006940.2| 149385 + tpg|BK006940.2| 148986 - INS 
 tpg|BK006941.2| 474327 + tpg|BK006941.2| 473692 - INS 
 tpg|BK006938.2| 1241105 + tpg|BK006938.2| 1241274 - INS 
 tpg|BK006940.2| 107964 + tpg|BK006940.2| 107256 - INS 
 tpg|BK006940.2| 64075 + tpg|BK006940.2| 64532 - INS 
 tpg|BK006940.2| 243253 + tpg|BK006940.2| 243113 - INS 
 tpg|BK006941.2| 987080 + tpg|BK006941.2| 986831 - INS 
 tpg|BK006940.2| 37194 + tpg|BK006940.2| 36583 - INS 
 tpg|BK006941.2| 744524 + tpg|BK006941.2| 744651 - INS 
 tpg|BK006940.2| 125610 + tpg|BK006940.2| 125284 - INS 
 tpg|BK006940.2| 240827 + tpg|BK006940.2| 240143 - INS 
 tpg|BK006938.2| 84113 + tpg|BK006938.2| 84869 - INS 
 tpg|BK006941.2| 355642 + tpg|BK006941.2| 355981 - INS 
 tpg|BK006940.2| 23229 + tpg|BK006940.2| 22761 - INS 
 tpg|BK006938.2| 1013121 + tpg|BK006938.2| 1013826 - INS 
 tpg|BK006940.2| 240192 + tpg|BK006940.2| 239564 - INS 
 tpg|BK006940.2| 251552 + tpg|BK006940.2| 251505 - INS 
 tpg|BK006941.2| 738888 + tpg|BK006941.2| 738288 - INS 
 tpg|BK006940.2| 32321 + tpg|BK006940.2| 31759 - INS 
 tpg|BK006941.2| 111772 + tpg|BK006941.2| 112021 - INS 
 tpg|BK006938.2| 1275311 + tpg|BK006938.2| 1275980 - INS 
 tpg|BK006940.2| 239334 + tpg|BK006940.2| 238923 - INS 
 tpg|BK006941.2| 465783 + tpg|BK006941.2| 465164 - INS 
 tpg|BK006940.2| 129695 + tpg|BK006940.2| 129010 - INS 
 tpg|BK006941.2| 108173 + tpg|BK006941.2| 107410 - INS 
 tpg|BK006938.2| 110925 + tpg|BK006938.2| 110181 - INS 
 tpg|BK006941.2| 765678 + tpg|BK006941.2| 766029 - INS 
 tpg|BK006938.2| 231221 + tpg|BK006938.2| 230891 - INS 
 tpg|BK006940.2| 115229 + tpg|BK006940.2| 115121 - INS 
 tpg|BK006941.2| 692430 + tpg|BK006941.2| 692335 - INS 
 tpg|BK006940.2| 214813 + tpg|BK006940.2| 215387 - INS 
 tpg|BK006938.2| 734577 + tpg|BK006938.2| 734433 - INS 
 tpg|BK006941.2| 130781 + tpg|BK006941.2| 130456 - INS 
 tpg|BK006941.2| 702192 + tpg|BK006941.2| 701808 - INS 
 tpg|BK006940.2| 55073 + tpg|BK006940.2| 55803 - INS 
 tpg|BK006940.2| 102195 + tpg|BK006940.2| 101493 - INS 
 tpg|BK006941.2| 205686 + tpg|BK006941.2| 205334 - INS 
 tpg|BK006941.2| 855132 + tpg|BK006941.2| 854430 - INS 
 tpg|BK006940.2| 228020 + tpg|BK006940.2| 228557 - INS 
 tpg|BK006941.2| 752234 + tpg|BK006941.2| 752415 - INS 
 tpg|BK006941.2| 758295 + tpg|BK006941.2| 758065 - INS 
 tpg|BK006940.2| 17213 + tpg|BK006940.2| 17072 - INS 
 tpg|BK006941.2| 797453 + tpg|BK006941.2| 796794 - INS 
 tpg|BK006938.2| 887108 + tpg|BK006938.2| 887674 - INS 
 tpg|BK006940.2| 146051 + tpg|BK006940.2| 145723 - INS 
 tpg|BK006941.2| 425802 + tpg|BK006941.2| 425201 - INS 
 tpg|BK006938.2| 124863 + tpg|BK006938.2| 124306 - INS 
 tpg|BK006940.2| 130939 + tpg|BK006940.2| 130534 - INS 
 tpg|BK006941.2| 831183 + tpg|BK006941.2| 830779 - INS 
 tpg|BK006941.2| 837607 + tpg|BK006941.2| 838357 - INS 
 tpg|BK006940.2| 176282 + tpg|BK006940.2| 176221 - INS 
 tpg|BK006941.2| 780706 + tpg|BK006941.2| 780817 - INS 
 tpg|BK006941.2| 920745 + tpg|BK006941.2| 920913 - INS 
 tpg|BK006941.2| 772183 + tpg|BK006941.2| 771410 - INS 
 tpg|BK006938.2| 267283 + tpg|BK006938.2| 267308 - INS 
 tpg|BK006941.2| 771458 + tpg|BK006941.2| 770881 - INS 
 tpg|BK006938.2| 207355 + tpg|BK006938.2| 207054 - INS 
 tpg|BK006941.2| 462541 + tpg|BK006941.2| 462166 - INS 
 tpg|BK006941.2| 754690 + tpg|BK006941.2| 754142 - INS 
 tpg|BK006938.2| 280101 + tpg|BK006938.2| 279489 - INS 
 tpg|BK006938.2| 1127795 + tpg|BK006938.2| 1127554 - INS 
 tpg|BK006941.2| 908358 + tpg|BK006941.2| 908057 - INS 
 tpg|BK006941.2| 56268 + tpg|BK006941.2| 55853 - INS 
 tpg|BK006938.2| 1420658 + tpg|BK006938.2| 1420364 - INS 
 tpg|BK006941.2| 245072 + tpg|BK006941.2| 244797 - INS 
 tpg|BK006941.2| 704359 + tpg|BK006941.2| 704101 - INS 
 tpg|BK006941.2| 700491 + tpg|BK006941.2| 699839 - INS 
 tpg|BK006941.2| 322632 + tpg|BK006941.2| 322108 - INS 
 tpg|BK006940.2| 108834 + tpg|BK006940.2| 108601 - INS 
 tpg|BK006941.2| 1014274 + tpg|BK006941.2| 1014240 - INS 
 tpg|BK006940.2| 39308 + tpg|BK006940.2| 38642 - INS 
 tpg|BK006941.2| 661456 + tpg|BK006941.2| 661801 - INS 
 tpg|BK006940.2| 14594 + tpg|BK006940.2| 14788 - INS 
 tpg|BK006941.2| 657339 + tpg|BK006941.2| 657673 - INS 
 tpg|BK006940.2| 177312 + tpg|BK006940.2| 177051 - INS 
 tpg|BK006941.2| 1019358 + tpg|BK006941.2| 1018833 - INS 
 tpg|BK006941.2| 651542 + tpg|BK006941.2| 650791 - INS 
 tpg|BK006940.2| 52977 + tpg|BK006940.2| 52848 - INS 
 tpg|BK006941.2| 311646 + tpg|BK006941.2| 311031 - INS 
 tpg|BK006938.2| 1395162 + tpg|BK006938.2| 1394922 - INS 
 tpg|BK006941.2| 1021869 + tpg|BK006941.2| 1021960 - INS 
 tpg|BK006940.2| 221512 + tpg|BK006940.2| 221527 - INS 
 tpg|BK006938.2| 395058 + tpg|BK006938.2| 394725 - INS 
 tpg|BK006940.2| 132738 + tpg|BK006940.2| 132770 - INS 
 tpg|BK006941.2| 639479 + tpg|BK006941.2| 638728 - INS 
 tpg|BK006940.2| 111889 + tpg|BK006940.2| 111686 - INS 
 tpg|BK006941.2| 1022907 + tpg|BK006941.2| 1022593 - INS 
 tpg|BK006940.2| 233651 + tpg|BK006940.2| 233604 - INS 
 tpg|BK006938.2| 1369497 + tpg|BK006938.2| 1369122 - INS 
 tpg|BK006940.2| 179132 + tpg|BK006940.2| 179275 - INS 
 tpg|BK006941.2| 1026519 + tpg|BK006941.2| 1026730 - INS 
 tpg|BK006940.2| 202991 + tpg|BK006940.2| 203467 - INS 
 tpg|BK006941.2| 10954 + tpg|BK006941.2| 11002 - INS 
 tpg|BK006938.2| 1299819 + tpg|BK006938.2| 1299576 - INS 
 tpg|BK006941.2| 13999 + tpg|BK006941.2| 14459 - INS 
 tpg|BK006940.2| 103883 + tpg|BK006940.2| 104459 - INS TTA
 tpg|BK006940.2| 219581 + tpg|BK006940.2| 219011 - INS 
 tpg|BK006941.2| 163637 + tpg|BK006941.2| 163264 - INS 
 tpg|BK006940.2| 248489 + tpg|BK006940.2| 247831 - INS 
 tpg|BK006941.2| 568379 + tpg|BK006941.2| 568359 - INS 
 tpg|BK006940.2| 51591 + tpg|BK006940.2| 51664 - INS GATA
 tpg|BK006940.2| 45060 + tpg|BK006940.2| 44447 - INS 
 tpg|BK006941.2| 554356 + tpg|BK006941.2| 554006 - INS 
 tpg|BK006941.2| 183492 + tpg|BK006941.2| 184072 - INS 
 tpg|BK006940.2| 15391 + tpg|BK006940.2| 15690 - INS 
 tpg|BK006938.2| 1351662 + tpg|BK006938.2| 1351487 - INS 
 tpg|BK006940.2| 163062 + tpg|BK006940.2| 162702 - INS 
 tpg|BK006941.2| 561796 + tpg|BK006941.2| 561704 - INS 
 tpg|BK006940.2| 56685 + tpg|BK006940.2| 56454 - INS 
 tpg|BK006940.2| 169809 + tpg|BK006940.2| 170088 - INS 
 tpg|BK006938.2| 484370 + tpg|BK006938.2| 484192 - INS 
 tpg|BK006941.2| 466967 + tpg|BK006941.2| 466202 - INS 
 tpg|BK006941.2| 857807 + tpg|BK006941.2| 857883 - INS 
 tpg|BK006940.2| 204461 + tpg|BK006940.2| 204090 - INS 
 tpg|BK006938.2| 1384121 + tpg|BK006938.2| 1384263 - INS 
 tpg|BK006938.2| 1252333 + tpg|BK006938.2| 1251637 - INS 
 tpg|BK006941.2| 207586 + tpg|BK006941.2| 208323 - INS 
 tpg|BK006940.2| 161736 + tpg|BK006940.2| 161288 - INS 
 tpg|BK006941.2| 904584 + tpg|BK006941.2| 904322 - INS 
 tpg|BK006940.2| 155986 + tpg|BK006940.2| 156470 - INS 
 tpg|BK006938.2| 1253438 + tpg|BK006938.2| 1252859 - INS 
 tpg|BK006941.2| 906366 + tpg|BK006941.2| 905887 - INS 
 tpg|BK006940.2| 256600 + tpg|BK006940.2| 257216 - INS 
 tpg|BK006940.2| 213288 + tpg|BK006940.2| 213009 - INS 
 tpg|BK006940.2| 152122 + tpg|BK006940.2| 152648 - INS 
 tpg|BK006938.2| 562647 + tpg|BK006938.2| 562086 - INS 
 tpg|BK006940.2| 19506 + tpg|BK006940.2| 18810 - INS 
 tpg|BK006941.2| 250510 + tpg|BK006941.2| 249832 - INS 
 tpg|BK006940.2| 6589 + tpg|BK006940.2| 6330 - INS 
 tpg|BK006940.2| 265495 + tpg|BK006940.2| 265834 - INS 
 tpg|BK006940.2| 73130 + tpg|BK006940.2| 72863 - INS 
 tpg|BK006940.2| 171169 + tpg|BK006940.2| 171377 - INS 
 tpg|BK006938.2| 601546 + tpg|BK006938.2| 601693 - INS 
 tpg|BK006941.2| 972193 + tpg|BK006941.2| 972271 - INS 
 tpg|BK006940.2| 267371 + tpg|BK006940.2| 267510 - INS 
 tpg|BK006940.2| 146774 + tpg|BK006940.2| 146351 - INS 
 tpg|BK006938.2| 398524 + tpg|BK006938.2| 398596 - INS 
 tpg|BK006940.2| 113575 + tpg|BK006940.2| 113572 - INS 
 tpg|BK006938.2| 366691 + tpg|BK006938.2| 367288 - INS 
 tpg|BK006940.2| 84752 + tpg|BK006940.2| 84389 - INS 
 tpg|BK006940.2| 231593 + tpg|BK006940.2| 231126 - INS 
 tpg|BK006938.2| 410196 + tpg|BK006938.2| 410868 - INS TCT
 tpg|BK006940.2| 268924 + tpg|BK006940.2| 268436 - INS 
 tpg|BK006941.2| 1006863 + tpg|BK006941.2| 1006405 - INS 
 tpg|BK006938.2| 88766 + tpg|BK006938.2| 88292 - INS 
 tpg|BK006941.2| 1007728 + tpg|BK006941.2| 1008232 - INS 
 tpg|BK006938.2| 927416 + tpg|BK006938.2| 927309 - INS 
 tpg|BK006941.2| 176032 + tpg|BK006941.2| 175531 - INS 
 tpg|BK006940.2| 262646 + tpg|BK006940.2| 262360 - INS 
 tpg|BK006938.2| 1378695 + tpg|BK006938.2| 1378629 - INS 
 tpg|BK006940.2| 90940 + tpg|BK006940.2| 90841 - INS 
 tpg|BK006941.2| 617418 + tpg|BK006941.2| 618073 - INS 
 tpg|BK006938.2| 479317 + tpg|BK006938.2| 479864 - INS 
 tpg|BK006940.2| 209165 + tpg|BK006940.2| 208577 - INS 
 tpg|BK006941.2| 40967 + tpg|BK006941.2| 40697 - INS 
 tpg|BK006940.2| 223681 + tpg|BK006940.2| 222944 - INS 
 tpg|BK006941.2| 689014 + tpg|BK006941.2| 689278 - INS 
 tpg|BK006940.2| 54407 + tpg|BK006940.2| 54127 - INS 
 tpg|BK006941.2| 868863 + tpg|BK006941.2| 869296 - INS 
 tpg|BK006940.2| 216348 + tpg|BK006940.2| 216305 - INS 
 tpg|BK006940.2| 209934 + tpg|BK006940.2| 210165 - INS 
 tpg|BK006941.2| 88432 + tpg|BK006941.2| 88350 - INS 
 tpg|BK006938.2| 477979 + tpg|BK006938.2| 477686 - INS 
 tpg|BK006940.2| 98436 + tpg|BK006940.2| 98516 - INS 
 tpg|BK006941.2| 86226 + tpg|BK006941.2| 86514 - INS 
 tpg|BK006940.2| 232508 + tpg|BK006940.2| 232395 - INS 
 tpg|BK006941.2| 91780 + tpg|BK006941.2| 91585 - INS 
 tpg|BK006940.2| 244812 + tpg|BK006940.2| 244764 - INS 
 tpg|BK006941.2| 826643 + tpg|BK006941.2| 826674 - INS 
 tpg|BK006938.2| 203791 + tpg|BK006938.2| 203534 - INS 
 tpg|BK006940.2| 39987 + tpg|BK006940.2| 40155 - INS 
 tpg|BK006941.2| 934217 + tpg|BK006941.2| 933868 - INS 
 tpg|BK006940.2| 166135 + tpg|BK006940.2| 166274 - INS 
 tpg|BK006941.2| 912050 + tpg|BK006941.2| 912102 - INS 
 tpg|BK006938.2| 444069 + tpg|BK006938.2| 444005 - INS 
 tpg|BK006941.2| 21016 + tpg|BK006941.2| 20819 - INS 
 tpg|BK006940.2| 196194 + tpg|BK006940.2| 195974 - INS 
 tpg|BK006938.2| 312532 + tpg|BK006938.2| 311801 - INS 
 tpg|BK006941.2| 825198 + tpg|BK006941.2| 824890 - INS 
 tpg|BK006940.2| 62452 + tpg|BK006940.2| 62801 - INS 
 tpg|BK006941.2| 168192 + tpg|BK006941.2| 167705 - INS 
 tpg|BK006941.2| 865793 + tpg|BK006941.2| 865156 - INS 
 tpg|BK006938.2| 343662 + tpg|BK006938.2| 343142 - INS 
 tpg|BK006940.2| 269511 + tpg|BK006940.2| 269159 - INS 
 tpg|BK006941.2| 37121 + tpg|BK006941.2| 36502 - INS 
 tpg|BK006938.2| 886544 + tpg|BK006938.2| 886237 - INS 
 tpg|BK006940.2| 68791 + tpg|BK006940.2| 69146 - INS 
 tpg|BK006941.2| 894548 + tpg|BK006941.2| 894051 - INS 
 tpg|BK006940.2| 95029 + tpg|BK006940.2| 95451 - INS 
 tpg|BK006938.2| 608930 + tpg|BK006938.2| 608998 - INS 
 tpg|BK006941.2| 431187 + tpg|BK006941.2| 430741 - INS 
 tpg|BK006941.2| 441681 + tpg|BK006941.2| 441291 - INS 
 tpg|BK006941.2| 472217 + tpg|BK006941.2| 472647 - INS 
 tpg|BK006940.2| 25457 + tpg|BK006940.2| 25017 - INS 
 tpg|BK006938.2| 1367147 + tpg|BK006938.2| 1367662 - INS 
 tpg|BK006941.2| 479781 + tpg|BK006941.2| 480271 - INS 
 tpg|BK006940.2| 118521 + tpg|BK006940.2| 118165 - INS 
 tpg|BK006938.2| 1250177 + tpg|BK006938.2| 1249609 - INS 
 tpg|BK006940.2| 48567 + tpg|BK006940.2| 48971 - INS 
 tpg|BK006941.2| 32206 + tpg|BK006941.2| 32165 - INS 
 tpg|BK006940.2| 229437 + tpg|BK006940.2| 229964 - INS 
 tpg|BK006940.2| 200345 + tpg|BK006940.2| 200239 - INS 
 tpg|BK006940.2| 255356 + tpg|BK006940.2| 255431 - INS 
 tpg|BK006941.2| 329468 + tpg|BK006941.2| 329228 - INS 
 tpg|BK006940.2| 88851 + tpg|BK006940.2| 88751 - INS 
 tpg|BK006941.2| 502639 + tpg|BK006941.2| 503225 - INS 
 tpg|BK006941.2| 691720 + tpg|BK006941.2| 691540 - INS 
 tpg|BK006940.2| 47684 + tpg|BK006940.2| 47425 - INS 
 tpg|BK006938.2| 210661 + tpg|BK006938.2| 210752 - INS 
 tpg|BK006940.2| 30335 + tpg|BK006940.2| 29943 - INS 
 tpg|BK006941.2| 320129 + tpg|BK006941.2| 320005 - INS 
 tpg|BK006940.2| 263785 + tpg|BK006940.2| 263955 - INS 
 tpg|BK006941.2| 22307 + tpg|BK006941.2| 22517 - INS 
 tpg|BK006940.2| 46404 + tpg|BK006940.2| 46171 - INS 
 tpg|BK006941.2| 316085 + tpg|BK006941.2| 315575 - INS 
 tpg|BK006940.2| 120211 + tpg|BK006940.2| 120597 - INS 
 tpg|BK006941.2| 653710 + tpg|BK006941.2| 654088 - INS 
 tpg|BK006938.2| 782042 + tpg|BK006938.2| 781835 - INS 
 tpg|BK006940.2| 74508 + tpg|BK006940.2| 74250 - INS 
 tpg|BK006941.2| 309729 + tpg|BK006941.2| 309683 - INS 
 tpg|BK006941.2| 532476 + tpg|BK006941.2| 532148 - INS 
 tpg|BK006940.2| 73753 + tpg|BK006940.2| 73695 - INS 
 tpg|BK006941.2| 595034 + tpg|BK006941.2| 595132 - INS 
 tpg|BK006940.2| 18553 + tpg|BK006940.2| 17857 - INS 
 tpg|BK006940.2| 172754 + tpg|BK006940.2| 172583 - INS 
 tpg|BK006938.2| 806085 + tpg|BK006938.2| 806650 - INS 
 tpg|BK006941.2| 281344 + tpg|BK006941.2| 281029 - INS 
 tpg|BK006940.2| 137363 + tpg|BK006940.2| 136961 - INS 
 tpg|BK006938.2| 746274 + tpg|BK006938.2| 746018 - INS 
 tpg|BK006940.2| 249404 + tpg|BK006940.2| 249371 - INS 
 tpg|BK006941.2| 585237 + tpg|BK006941.2| 584488 - INS 
 tpg|BK006940.2| 150362 + tpg|BK006940.2| 150089 - INS 
 tpg|BK006940.2| 129125 + tpg|BK006940.2| 128440 - INS 
 tpg|BK006938.2| 103562 + tpg|BK006938.2| 102864 - INS 
 tpg|BK006941.2| 555042 + tpg|BK006941.2| 554616 - INS 
 tpg|BK006940.2| 41125 + tpg|BK006940.2| 40952 - INS 
 tpg|BK006941.2| 159689 + tpg|BK006941.2| 160170 - INS 
 tpg|BK006941.2| 1041846 + tpg|BK006941.2| 1042584 - INS 
 tpg|BK006941.2| 1008795 + tpg|BK006941.2| 1009337 - INS 
 tpg|BK006940.2| 188251 + tpg|BK006940.2| 188463 - INS 
 tpg|BK006940.2| 66428 + tpg|BK006940.2| 66272 - INS 
 tpg|BK006941.2| 680601 + tpg|BK006941.2| 680177 - INS 
 tpg|BK006940.2| 85292 + tpg|BK006940.2| 85505 - INS 
 tpg|BK006941.2| 332845 + tpg|BK006941.2| 333043 - INS 
 tpg|BK006940.2| 144703 + tpg|BK006940.2| 144792 - INS 
 tpg|BK006940.2| 121589 + tpg|BK006940.2| 122333 - INS 
 tpg|BK006941.2| 715055 + tpg|BK006941.2| 715735 - INS 
 tpg|BK006940.2| 180089 + tpg|BK006940.2| 179777 - INS 
 tpg|BK006941.2| 721686 + tpg|BK006941.2| 722212 - INS 
 tpg|BK006941.2| 486117 + tpg|BK006941.2| 485398 - INS 
 tpg|BK006940.2| 70058 + tpg|BK006940.2| 69868 - INS 
 tpg|BK006941.2| 681199 + tpg|BK006941.2| 680752 - INS 
 tpg|BK006940.2| 35489 + tpg|BK006940.2| 36126 - INS 
 tpg|BK006940.2| 61118 + tpg|BK006940.2| 61006 - INS 
 tpg|BK006941.2| 1045593 + tpg|BK006941.2| 1045386 - INS 
 tpg|BK006940.2| 34935 + tpg|BK006940.2| 34330 - INS 
 tpg|BK006941.2| 549537 + tpg|BK006941.2| 549157 - INS 
 tpg|BK006941.2| 674055 + tpg|BK006941.2| 673859 - INS 
 tpg|BK006940.2| 241325 + tpg|BK006940.2| 240832 - INS 
 tpg|BK006941.2| 209300 + tpg|BK006941.2| 209435 - INS 
 tpg|BK006940.2| 178112 + tpg|BK006940.2| 177691 - INS 
 tpg|BK006938.2| 1478330 + tpg|BK006938.2| 1477891 - INS 
 tpg|BK006940.2| 102796 + tpg|BK006940.2| 102250 - INS 
 tpg|BK006941.2| 451282 + tpg|BK006941.2| 450695 - INS 
 tpg|BK006940.2| 173458 + tpg|BK006940.2| 173336 - INS 
 tpg|BK006941.2| 496384 + tpg|BK006941.2| 496024 - INS 
 tpg|BK006938.2| 643977 + tpg|BK006938.2| 643210 - INS 
 tpg|BK006940.2| 59332 + tpg|BK006940.2| 59500 - INS 
 tpg|BK006941.2| 696268 + tpg|BK006941.2| 696528 - INS 
 tpg|BK006941.2| 713807 + tpg|BK006941.2| 713896 - INS 
 tpg|BK006941.2| 726121 + tpg|BK006941.2| 725761 - INS 
 tpg|BK006938.2| 620174 + tpg|BK006938.2| 619981 - INS 
 tpg|BK006941.2| 117395 + tpg|BK006941.2| 117985 - INS 
 tpg|BK006938.2| 625853 + tpg|BK006938.2| 625399 - INS 
 tpg|BK006941.2| 836681 + tpg|BK006941.2| 836844 - INS 
 tpg|BK006941.2| 399519 + tpg|BK006941.2| 399948 - INS 
 tpg|BK006941.2| 19372 + tpg|BK006941.2| 19984 - INS 
 tpg|BK006941.2| 807433 + tpg|BK006941.2| 808007 - INS 
 tpg|BK006938.2| 1002003 + tpg|BK006938.2| 1002266 - INS 
 tpg|BK006941.2| 161065 + tpg|BK006941.2| 160680 - INS 
 tpg|BK006941.2| 608957 + tpg|BK006941.2| 609276 - INS 
 tpg|BK006938.2| 1020959 + tpg|BK006938.2| 1020579 - INS 
 tpg|BK006940.2| 112809 + tpg|BK006940.2| 112658 - INS 
 tpg|BK006941.2| 142115 + tpg|BK006941.2| 141512 - INS 
 tpg|BK006940.2| 245844 + tpg|BK006940.2| 245379 - INS 
 tpg|BK006940.2| 153652 + tpg|BK006940.2| 153369 - INS 
 tpg|BK006940.2| 234771 + tpg|BK006940.2| 234363 - INS 
 tpg|BK006941.2| 71610 + tpg|BK006941.2| 71263 - INS 
 tpg|BK006940.2| 235626 + tpg|BK006940.2| 236069 - INS 
 tpg|BK006938.2| 1057874 + tpg|BK006938.2| 1057739 - INS 
 tpg|BK006940.2| 264461 + tpg|BK006940.2| 264624 - INS 
 tpg|BK006940.2| 266851 + tpg|BK006940.2| 266474 - INS 
 tpg|BK006940.2| 131799 + tpg|BK006940.2| 131957 - INS 
 tpg|BK006941.2| 434867 + tpg|BK006941.2| 434719 - INS 
 tpg|BK006940.2| 62004 + tpg|BK006940.2| 61372 - INS 
 tpg|BK006938.2| 569621 + tpg|BK006938.2| 569896 - INS 
 tpg|BK006940.2| 32755 + tpg|BK006940.2| 32561 - INS 
 tpg|BK006941.2| 755134 + tpg|BK006941.2| 754899 - INS 
 tpg|BK006940.2| 8958 + tpg|BK006940.2| 8624 - INS 
 tpg|BK006941.2| 202832 + tpg|BK006941.2| 203283 - INS 
 tpg|BK006940.2| 86585 + tpg|BK006940.2| 86358 - INS 
 tpg|BK006938.2| 566239 + tpg|BK006938.2| 565654 - INS 
 tpg|BK006940.2| 160591 + tpg|BK006940.2| 160358 - INS 
 tpg|BK006941.2| 217288 + tpg|BK006941.2| 217809 - INS 
 tpg|BK006940.2| 137922 + tpg|BK006940.2| 137566 - INS 
 tpg|BK006941.2| 169029 + tpg|BK006941.2| 168328 - INS 
 tpg|BK006940.2| 13463 + tpg|BK006940.2| 13310 - INS 
 tpg|BK006938.2| 924386 + tpg|BK006938.2| 924560 - INS 
 tpg|BK006940.2| 186541 + tpg|BK006940.2| 187290 - INS 
 tpg|BK006941.2| 164911 + tpg|BK006941.2| 165657 - INS 
 tpg|BK006940.2| 25834 + tpg|BK006940.2| 26003 - INS 
 tpg|BK006940.2| 207000 + tpg|BK006940.2| 206597 - INS 
 tpg|BK006938.2| 164079 + tpg|BK006938.2| 163992 - INS 
 tpg|BK006940.2| 97279 + tpg|BK006940.2| 97235 - INS 
 tpg|BK006940.2| 201019 + tpg|BK006940.2| 201081 - INS 
 tpg|BK006940.2| 238075 + tpg|BK006940.2| 237722 - INS 
 tpg|BK006938.2| 314331 + tpg|BK006938.2| 313966 - INS 
 tpg|BK006941.2| 889611 + tpg|BK006941.2| 888844 - INS 
 tpg|BK006941.2| 219239 + tpg|BK006941.2| 219034 - INS 
 tpg|BK006938.2| 1217408 + tpg|BK006938.2| 1216843 - INS 
 tpg|BK006941.2| 392558 + tpg|BK006941.2| 393237 - INS 
 tpg|BK006941.2| 895271 + tpg|BK006941.2| 895204 - INS 
 tpg|BK006941.2| 235702 + tpg|BK006941.2| 235965 - INS 
 tpg|BK006938.2| 176472 + tpg|BK006938.2| 176460 - INS 
 tpg|BK006941.2| 366047 + tpg|BK006941.2| 365808 - INS 
 tpg|BK006941.2| 462977 + tpg|BK006941.2| 463251 - INS 
 tpg|BK006938.2| 177814 + tpg|BK006938.2| 177523 - INS 
 tpg|BK006941.2| 947444 + tpg|BK006941.2| 946953 - INS 
 tpg|BK006941.2| 966350 + tpg|BK006941.2| 966184 - INS 
 tpg|BK006938.2| 977156 + tpg|BK006938.2| 977335 - INS 
 tpg|BK006941.2| 970482 + tpg|BK006941.2| 970243 - INS 
 tpg|BK006938.2| 1164151 + tpg|BK006938.2| 1164629 - INS 
 tpg|BK006941.2| 251097 + tpg|BK006941.2| 251530 - INS 
 tpg|BK006941.2| 122556 + tpg|BK006941.2| 121792 - INS 
 tpg|BK006938.2| 1445303 + tpg|BK006938.2| 1445366 - INS 
 tpg|BK006941.2| 498496 + tpg|BK006941.2| 498157 - INS 
 tpg|BK006941.2| 29540 + tpg|BK006941.2| 29793 - INS 
 tpg|BK006938.2| 373546 + tpg|BK006938.2| 373896 - INS 
 tpg|BK006941.2| 1000895 + tpg|BK006941.2| 1001351 - INS 
 tpg|BK006941.2| 326279 + tpg|BK006941.2| 325935 - INS 
 tpg|BK006938.2| 292644 + tpg|BK006938.2| 292972 - INS 
 tpg|BK006941.2| 1025650 + tpg|BK006941.2| 1024907 - INS 
 tpg|BK006941.2| 551844 + tpg|BK006941.2| 552073 - INS 
 tpg|BK006941.2| 1048545 + tpg|BK006941.2| 1048124 - INS 
 tpg|BK006938.2| 1141773 + tpg|BK006938.2| 1141676 - INS 
 tpg|BK006941.2| 1076462 + tpg|BK006941.2| 1075706 - INS 
 tpg|BK006941.2| 836086 + tpg|BK006941.2| 835864 - INS 
 tpg|BK006938.2| 87413 + tpg|BK006938.2| 87397 - INS 
 tpg|BK006938.2| 342250 + tpg|BK006938.2| 342686 - INS 
 tpg|BK006938.2| 786863 + tpg|BK006938.2| 787271 - INS 
 tpg|BK006938.2| 22032 + tpg|BK006938.2| 22281 - INS 
 tpg|BK006938.2| 857805 + tpg|BK006938.2| 858307 - INS 
 tpg|BK006941.2| 106364 + tpg|BK006941.2| 105680 - INS 
 tpg|BK006941.2| 99188 + tpg|BK006941.2| 99963 - INS 
 tpg|BK006941.2| 456251 + tpg|BK006941.2| 456914 - INS 
 tpg|BK006941.2| 775881 + tpg|BK006941.2| 776457 - INS 
 tpg|BK006941.2| 802689 + tpg|BK006941.2| 803003 - INS 
 tpg|BK006941.2| 95045 + tpg|BK006941.2| 95349 - INS 
 tpg|BK006941.2| 896942 + tpg|BK006941.2| 896490 - INS 
 tpg|BK006941.2| 477896 + tpg|BK006941.2| 477603 - INS 
 tpg|BK006941.2| 159063 + tpg|BK006941.2| 158439 - INS 
 tpg|BK006938.2| 1347552 + tpg|BK006938.2| 1347660 - INS 
 tpg|BK006938.2| 56228 + tpg|BK006938.2| 56360 - INS 
 tpg|BK006938.2| 37518 + tpg|BK006938.2| 37757 - INS 
 tpg|BK006941.2| 228596 + tpg|BK006941.2| 228144 - INS 
 tpg|BK006941.2| 194566 + tpg|BK006941.2| 194551 - INS 
 tpg|BK006938.2| 237849 + tpg|BK006938.2| 238428 - INS 
 tpg|BK006938.2| 420661 + tpg|BK006938.2| 420496 - INS 
 tpg|BK006941.2| 628929 + tpg|BK006941.2| 629366 - INS 
 tpg|BK006938.2| 1310461 + tpg|BK006938.2| 1311202 - INS 
 tpg|BK006938.2| 1284564 + tpg|BK006938.2| 1284009 - INS 
 tpg|BK006941.2| 275887 + tpg|BK006941.2| 275313 - INS 
 tpg|BK006938.2| 754064 + tpg|BK006938.2| 754105 - INS 
 tpg|BK006941.2| 1066107 + tpg|BK006941.2| 1066180 - INS 
 tpg|BK006941.2| 238430 + tpg|BK006941.2| 238730 - INS 
 tpg|BK006938.2| 315379 + tpg|BK006938.2| 315592 - INS 
 tpg|BK006941.2| 274781 + tpg|BK006941.2| 274404 - INS 
 tpg|BK006941.2| 1003350 + tpg|BK006941.2| 1003169 - INS 
 tpg|BK006941.2| 919625 + tpg|BK006941.2| 920042 - INS 
 tpg|BK006938.2| 473150 + tpg|BK006938.2| 473398 - INS 
 tpg|BK006941.2| 917483 + tpg|BK006941.2| 918140 - INS 
 tpg|BK006938.2| 1157263 + tpg|BK006938.2| 1156530 - INS 
 tpg|BK006938.2| 1144087 + tpg|BK006938.2| 1143336 - INS 
 tpg|BK006941.2| 234954 + tpg|BK006941.2| 234608 - INS 
 tpg|BK006938.2| 500152 + tpg|BK006938.2| 499715 - INS 
 tpg|BK006941.2| 637441 + tpg|BK006941.2| 637683 - INS 
 tpg|BK006941.2| 289258 + tpg|BK006941.2| 289442 - INS 
 tpg|BK006941.2| 385556 + tpg|BK006941.2| 385957 - INS 
 tpg|BK006941.2| 519859 + tpg|BK006941.2| 520363 - INS 
 tpg|BK006941.2| 517152 + tpg|BK006941.2| 516501 - INS 
 tpg|BK006941.2| 504832 + tpg|BK006941.2| 504681 - INS 
 tpg|BK006938.2| 1385913 + tpg|BK006938.2| 1385571 - INS 
 tpg|BK006941.2| 137563 + tpg|BK006941.2| 137471 - INS 
 tpg|BK006941.2| 335242 + tpg|BK006941.2| 335176 - INS 
 tpg|BK006938.2| 363768 + tpg|BK006938.2| 363675 - INS 
 tpg|BK006941.2| 973420 + tpg|BK006941.2| 973946 - INS 
 tpg|BK006941.2| 252028 + tpg|BK006941.2| 252052 - INS 
 tpg|BK006938.2| 945468 + tpg|BK006938.2| 944957 - INS 
 tpg|BK006941.2| 843719 + tpg|BK006941.2| 843855 - INS 
 tpg|BK006938.2| 967259 + tpg|BK006938.2| 966510 - INS 
 tpg|BK006941.2| 727344 + tpg|BK006941.2| 728095 - INS 
 tpg|BK006941.2| 45261 + tpg|BK006941.2| 45332 - INS 
 tpg|BK006938.2| 558111 + tpg|BK006938.2| 557450 - INS 
 tpg|BK006941.2| 295953 + tpg|BK006941.2| 295443 - INS 
 tpg|BK006941.2| 767505 + tpg|BK006941.2| 767822 - INS 
 tpg|BK006938.2| 1435408 + tpg|BK006938.2| 1435054 - INS 
 tpg|BK006941.2| 366632 + tpg|BK006941.2| 367141 - INS 
 tpg|BK006941.2| 48312 + tpg|BK006941.2| 47667 - INS 
 tpg|BK006938.2| 1063703 + tpg|BK006938.2| 1063136 - INS 
 tpg|BK006941.2| 939979 + tpg|BK006941.2| 939733 - INS 
 tpg|BK006941.2| 932762 + tpg|BK006941.2| 932373 - INS 
 tpg|BK006938.2| 612948 + tpg|BK006938.2| 612723 - INS 
 tpg|BK006941.2| 884267 + tpg|BK006941.2| 884023 - INS 
 tpg|BK006938.2| 261772 + tpg|BK006938.2| 261287 - INS 
 tpg|BK006941.2| 522068 + tpg|BK006941.2| 521694 - INS 
 tpg|BK006938.2| 1328044 + tpg|BK006938.2| 1327698 - INS 
 tpg|BK006941.2| 92505 + tpg|BK006941.2| 92180 - INS 
 tpg|BK006941.2| 681643 + tpg|BK006941.2| 682355 - INS 
 tpg|BK006941.2| 491693 + tpg|BK006941.2| 492143 - INS 
 tpg|BK006941.2| 206837 + tpg|BK006941.2| 207071 - INS 
 tpg|BK006941.2| 1080774 + tpg|BK006941.2| 1081053 - INS 
 tpg|BK006938.2| 1259050 + tpg|BK006938.2| 1258768 - INS 
 tpg|BK006941.2| 850536 + tpg|BK006941.2| 851101 - INS 
 tpg|BK006941.2| 908908 + tpg|BK006941.2| 908819 - INS 
 tpg|BK006938.2| 712276 + tpg|BK006938.2| 711914 - INS 
 tpg|BK006941.2| 270221 + tpg|BK006941.2| 270844 - INS 
 tpg|BK006941.2| 1017187 + tpg|BK006941.2| 1016501 - INS 
 tpg|BK006941.2| 1036095 + tpg|BK006941.2| 1035442 - INS 
 tpg|BK006941.2| 155908 + tpg|BK006941.2| 155532 - INS 
 tpg|BK006941.2| 785261 + tpg|BK006941.2| 784794 - INS 
 tpg|BK006938.2| 1518975 + tpg|BK006938.2| 1519208 - INS 
 tpg|BK006938.2| 833996 + tpg|BK006938.2| 833697 - INS 
 tpg|BK006938.2| 838718 + tpg|BK006938.2| 839200 - INS 
 tpg|BK006938.2| 718080 + tpg|BK006938.2| 718625 - INS 
 tpg|BK006938.2| 106977 + tpg|BK006938.2| 106681 - INS 
 tpg|BK006938.2| 683169 + tpg|BK006938.2| 682756 - INS 
 tpg|BK006938.2| 638925 + tpg|BK006938.2| 638580 - INS 
 tpg|BK006938.2| 617554 + tpg|BK006938.2| 617066 - INS 
 tpg|BK006941.2| 83043 + tpg|BK006941.2| 83249 - INS 
 tpg|BK006938.2| 1045155 + tpg|BK006938.2| 1045076 - INS 
 tpg|BK006938.2| 1415623 + tpg|BK006938.2| 1415111 - INS 
 tpg|BK006938.2| 1087847 + tpg|BK006938.2| 1088367 - INS 
 tpg|BK006938.2| 502459 + tpg|BK006938.2| 502293 - INS 
 tpg|BK006941.2| 905775 + tpg|BK006941.2| 905052 - INS 
 tpg|BK006941.2| 890756 + tpg|BK006941.2| 890805 - INS 
 tpg|BK006938.2| 474419 + tpg|BK006938.2| 473879 - INS 
 tpg|BK006941.2| 881739 + tpg|BK006941.2| 881615 - INS 
 tpg|BK006941.2| 386993 + tpg|BK006941.2| 386743 - INS 
 tpg|BK006941.2| 847739 + tpg|BK006941.2| 847990 - INS 
 tpg|BK006941.2| 364416 + tpg|BK006941.2| 364021 - INS 
 tpg|BK006938.2| 1158352 + tpg|BK006938.2| 1158244 - INS 
 tpg|BK006941.2| 361663 + tpg|BK006941.2| 361567 - INS 
 tpg|BK006941.2| 960212 + tpg|BK006941.2| 959634 - INS 
 tpg|BK006941.2| 202263 + tpg|BK006941.2| 202154 - INS 
 tpg|BK006938.2| 1391963 + tpg|BK006938.2| 1391655 - INS 
 tpg|BK006941.2| 253411 + tpg|BK006941.2| 252669 - INS 
 tpg|BK006941.2| 705530 + tpg|BK006941.2| 705326 - INS 
 tpg|BK006938.2| 423598 + tpg|BK006938.2| 423199 - INS 
 tpg|BK006941.2| 683446 + tpg|BK006941.2| 683622 - INS 
 tpg|BK006938.2| 1248807 + tpg|BK006938.2| 1248943 - INS 
 tpg|BK006941.2| 852540 + tpg|BK006941.2| 852999 - INS 
 tpg|BK006941.2| 517941 + tpg|BK006941.2| 517776 - INS 
 tpg|BK006941.2| 1020859 + tpg|BK006941.2| 1020338 - INS 
 tpg|BK006941.2| 639935 + tpg|BK006941.2| 639227 - INS 
 tpg|BK006941.2| 308422 + tpg|BK006941.2| 308278 - INS 
 tpg|BK006941.2| 150520 + tpg|BK006941.2| 151075 - INS 
 tpg|BK006941.2| 788025 + tpg|BK006941.2| 787910 - INS 
 tpg|BK006941.2| 900452 + tpg|BK006941.2| 900377 - INS 
 tpg|BK006941.2| 604258 + tpg|BK006941.2| 603786 - INS 
 tpg|BK006941.2| 596193 + tpg|BK006941.2| 596097 - INS 
 tpg|BK006938.2| 217474 + tpg|BK006938.2| 217166 - INS 
 tpg|BK006941.2| 25104 + tpg|BK006941.2| 25610 - INS 
 tpg|BK006941.2| 1073372 + tpg|BK006941.2| 1073988 - INS 
 tpg|BK006941.2| 427914 + tpg|BK006941.2| 427339 - INS 
 tpg|BK006941.2| 1079598 + tpg|BK006941.2| 1079523 - INS 
 tpg|BK006941.2| 610064 + tpg|BK006941.2| 609947 - INS 
 tpg|BK006941.2| 44591 + tpg|BK006941.2| 44190 - INS 
 tpg|BK006941.2| 283628 + tpg|BK006941.2| 284119 - INS 
 tpg|BK006938.2| 1485617 + tpg|BK006938.2| 1485232 - INS 
 tpg|BK006941.2| 916572 + tpg|BK006941.2| 916638 - INS 
 tpg|BK006938.2| 60035 + tpg|BK006938.2| 59972 - INS 
 tpg|BK006941.2| 152517 + tpg|BK006941.2| 152500 - INS 
 tpg|BK006941.2| 43905 + tpg|BK006941.2| 43403 - INS 
 tpg|BK006941.2| 635521 + tpg|BK006941.2| 635046 - INS 
 tpg|BK006938.2| 1170690 + tpg|BK006938.2| 1170600 - INS 
 tpg|BK006941.2| 717811 + tpg|BK006941.2| 718040 - INS 
 tpg|BK006941.2| 64642 + tpg|BK006941.2| 64588 - INS 
 tpg|BK006938.2| 731824 + tpg|BK006938.2| 731361 - INS 
 tpg|BK006938.2| 125979 + tpg|BK006938.2| 125898 - INS 
 tpg|BK006941.2| 876492 + tpg|BK006941.2| 875802 - INS 
 tpg|BK006938.2| 947064 + tpg|BK006938.2| 947210 - INS 
 tpg|BK006938.2| 637082 + tpg|BK006938.2| 637052 - INS 
 tpg|BK006941.2| 215978 + tpg|BK006941.2| 215599 - INS 
 tpg|BK006938.2| 1146928 + tpg|BK006938.2| 1146910 - INS 
 tpg|BK006938.2| 1137030 + tpg|BK006938.2| 1136992 - INS 
 tpg|BK006941.2| 791009 + tpg|BK006941.2| 790606 - INS 
 tpg|BK006941.2| 457892 + tpg|BK006941.2| 457819 - INS 
 tpg|BK006938.2| 1328631 + tpg|BK006938.2| 1329361 - INS 
 tpg|BK006941.2| 212763 + tpg|BK006941.2| 212600 - INS 
 tpg|BK006941.2| 903468 + tpg|BK006941.2| 903843 - INS 
 tpg|BK006941.2| 442170 + tpg|BK006941.2| 442664 - INS 
 tpg|BK006938.2| 1428730 + tpg|BK006938.2| 1428673 - INS 
 tpg|BK006941.2| 1063855 + tpg|BK006941.2| 1064142 - INS 
 tpg|BK006938.2| 571318 + tpg|BK006938.2| 570789 - INS 
 tpg|BK006941.2| 809953 + tpg|BK006941.2| 809371 - INS 
 tpg|BK006941.2| 832070 + tpg|BK006941.2| 832562 - INS 
 tpg|BK006941.2| 490378 + tpg|BK006941.2| 489732 - INS 
 tpg|BK006938.2| 1338442 + tpg|BK006938.2| 1338467 - INS 
 tpg|BK006938.2| 848829 + tpg|BK006938.2| 848839 - INS 
 tpg|BK006941.2| 296573 + tpg|BK006941.2| 296063 - INS 
 tpg|BK006941.2| 188918 + tpg|BK006941.2| 188577 - INS 
 tpg|BK006941.2| 1055999 + tpg|BK006941.2| 1055629 - INS 
 tpg|BK006938.2| 1357388 + tpg|BK006938.2| 1357124 - INS 
 tpg|BK006941.2| 18626 + tpg|BK006941.2| 17918 - INS 
 tpg|BK006941.2| 673547 + tpg|BK006941.2| 673004 - INS 
 tpg|BK006938.2| 509126 + tpg|BK006938.2| 508406 - INS 
 tpg|BK006941.2| 936515 + tpg|BK006941.2| 937041 - INS 
 tpg|BK006938.2| 96110 + tpg|BK006938.2| 96702 - INS 
 tpg|BK006938.2| 1238058 + tpg|BK006938.2| 1237397 - INS 
 tpg|BK006941.2| 437111 + tpg|BK006941.2| 437481 - INS 
 tpg|BK006938.2| 168733 + tpg|BK006938.2| 169452 - INS 
 tpg|BK006941.2| 182449 + tpg|BK006941.2| 183118 - INS 
 tpg|BK006941.2| 146221 + tpg|BK006941.2| 146585 - INS 
 tpg|BK006941.2| 172682 + tpg|BK006941.2| 173078 - INS 
 tpg|BK006938.2| 976020 + tpg|BK006938.2| 976413 - INS 
 tpg|BK006938.2| 439860 + tpg|BK006938.2| 440248 - INS 
 tpg|BK006941.2| 888009 + tpg|BK006941.2| 887610 - INS 
 tpg|BK006941.2| 288530 + tpg|BK006941.2| 288342 - INS 
 tpg|BK006941.2| 795378 + tpg|BK006941.2| 795181 - INS 
 tpg|BK006938.2| 1449903 + tpg|BK006938.2| 1449613 - INS 
 tpg|BK006941.2| 611366 + tpg|BK006941.2| 610663 - INS 
 tpg|BK006941.2| 485337 + tpg|BK006941.2| 484992 - INS 
 tpg|BK006941.2| 354037 + tpg|BK006941.2| 353542 - INS 
 tpg|BK006938.2| 793504 + tpg|BK006938.2| 793224 - INS 
 tpg|BK006941.2| 458623 + tpg|BK006941.2| 458299 - INS 
 tpg|BK006941.2| 455148 + tpg|BK006941.2| 455121 - INS 
 tpg|BK006938.2| 1355294 + tpg|BK006938.2| 1354738 - INS 
 tpg|BK006941.2| 141484 + tpg|BK006941.2| 140922 - INS 
 tpg|BK006941.2| 825721 + tpg|BK006941.2| 825567 - INS 
 tpg|BK006941.2| 306127 + tpg|BK006941.2| 306712 - INS 
 tpg|BK006938.2| 1073604 + tpg|BK006938.2| 1073012 - INS 
 tpg|BK006941.2| 254005 + tpg|BK006941.2| 253504 - INS 
 tpg|BK006938.2| 195198 + tpg|BK006938.2| 195836 - INS 
 tpg|BK006941.2| 525751 + tpg|BK006941.2| 525197 - INS 
 tpg|BK006938.2| 1294254 + tpg|BK006938.2| 1293938 - INS 
 tpg|BK006941.2| 459298 + tpg|BK006941.2| 458801 - INS 
 tpg|BK006941.2| 69891 + tpg|BK006941.2| 69758 - INS 
 tpg|BK006941.2| 944449 + tpg|BK006941.2| 944344 - INS 
 tpg|BK006941.2| 369362 + tpg|BK006941.2| 368618 - INS 
 tpg|BK006938.2| 252682 + tpg|BK006938.2| 252880 - INS 
 tpg|BK006941.2| 954308 + tpg|BK006941.2| 954290 - INS 
 tpg|BK006938.2| 242513 + tpg|BK006938.2| 241748 - INS 
 tpg|BK006938.2| 1496727 + tpg|BK006938.2| 1496779 - INS 
 tpg|BK006941.2| 374872 + tpg|BK006941.2| 374837 - INS 
 tpg|BK006941.2| 560843 + tpg|BK006941.2| 560581 - INS 
 tpg|BK006941.2| 764148 + tpg|BK006941.2| 763710 - INS 
 tpg|BK006941.2| 914742 + tpg|BK006941.2| 914902 - INS 
 tpg|BK006941.2| 896284 + tpg|BK006941.2| 895756 - INS 
 tpg|BK006941.2| 955149 + tpg|BK006941.2| 954658 - INS 
 tpg|BK006938.2| 636348 + tpg|BK006938.2| 636272 - INS 
 tpg|BK006941.2| 388477 + tpg|BK006941.2| 388035 - INS 
 tpg|BK006941.2| 897599 + tpg|BK006941.2| 897745 - INS 
 tpg|BK006938.2| 689080 + tpg|BK006938.2| 688464 - INS 
 tpg|BK006941.2| 862263 + tpg|BK006941.2| 862588 - INS 
 tpg|BK006938.2| 755877 + tpg|BK006938.2| 755260 - INS 
 tpg|BK006941.2| 436337 + tpg|BK006941.2| 435616 - INS  tpg|BK006938.2| 
 tpg|BK006941.2| 436337 + tpg|BK006941.2| 435616 - INS  tpg|BK006938.2| 
556172 + tpg|BK006938.2| 556556 - INS 
 tpg|BK006941.2| 3884 + tpg|BK006941.2| 3426 - INS 
 tpg|BK006941.2| 765230 + tpg|BK006941.2| 764959 - INS 
 tpg|BK006941.2| 694356 + tpg|BK006941.2| 694222 - INS 
 tpg|BK006941.2| 482369 + tpg|BK006941.2| 481988 - INS 
 tpg|BK006938.2| 1107294 + tpg|BK006938.2| 1106520 - INS 
 tpg|BK006941.2| 397024 + tpg|BK006941.2| 397422 - INS 
 tpg|BK006938.2| 288577 + tpg|BK006938.2| 288982 - INS 
 tpg|BK006941.2| 953449 + tpg|BK006941.2| 953309 - INS 
 tpg|BK006938.2| 300048 + tpg|BK006938.2| 299660 - INS 
 tpg|BK006941.2| 943891 + tpg|BK006941.2| 943443 - INS 
 tpg|BK006941.2| 108504 + tpg|BK006941.2| 108161 - INS 
 tpg|BK006938.2| 26584 + tpg|BK006938.2| 26123 - INS 
 tpg|BK006941.2| 994014 + tpg|BK006941.2| 993442 - INS 
 tpg|BK006941.2| 254662 + tpg|BK006941.2| 254273 - INS 
 tpg|BK006938.2| 977646 + tpg|BK006938.2| 978280 - INS 
 tpg|BK006941.2| 324872 + tpg|BK006941.2| 324586 - INS 
 tpg|BK006941.2| 255438 + tpg|BK006941.2| 256065 - INS 
 tpg|BK006941.2| 1029707 + tpg|BK006941.2| 1030246 - INS A
 tpg|BK006941.2| 186470 + tpg|BK006941.2| 186360 - INS 
 tpg|BK006941.2| 231356 + tpg|BK006941.2| 230728 - INS 
 tpg|BK006941.2| 512629 + tpg|BK006941.2| 512128 - INS 
 tpg|BK006938.2| 1194376 + tpg|BK006938.2| 1194500 - INS 
 tpg|BK006941.2| 675456 + tpg|BK006941.2| 675099 - INS 
 tpg|BK006941.2| 323806 + tpg|BK006941.2| 323373 - INS 
 tpg|BK006938.2| 962813 + tpg|BK006938.2| 962630 - INS 
 tpg|BK006938.2| 542513 + tpg|BK006938.2| 543056 - INS 
 tpg|BK006941.2| 312221 + tpg|BK006941.2| 312650 - INS 
 tpg|BK006941.2| 93031 + tpg|BK006941.2| 92820 - INS 
 tpg|BK006938.2| 1272359 + tpg|BK006938.2| 1271736 - INS 
 tpg|BK006941.2| 300676 + tpg|BK006941.2| 300226 - INS 
 tpg|BK006938.2| 225780 + tpg|BK006938.2| 225630 - INS 
 tpg|BK006941.2| 469292 + tpg|BK006941.2| 468708 - INS 
 tpg|BK006941.2| 419773 + tpg|BK006941.2| 419801 - INS 
 tpg|BK006938.2| 709073 + tpg|BK006938.2| 708790 - INS 
 tpg|BK006938.2| 215861 + tpg|BK006938.2| 215266 - INS 
 tpg|BK006938.2| 700405 + tpg|BK006938.2| 700550 - INS 
 tpg|BK006941.2| 171806 + tpg|BK006941.2| 171555 - INS 
 tpg|BK006941.2| 72063 + tpg|BK006941.2| 72083 - INS 
 tpg|BK006938.2| 848145 + tpg|BK006938.2| 847451 - INS 
 tpg|BK006941.2| 644522 + tpg|BK006941.2| 644025 - INS 
 tpg|BK006941.2| 263526 + tpg|BK006941.2| 262948 - INS 
 tpg|BK006941.2| 628567 + tpg|BK006941.2| 628394 - INS 
 tpg|BK006938.2| 1213837 + tpg|BK006938.2| 1213523 - INS 
 tpg|BK006941.2| 742045 + tpg|BK006941.2| 742181 - INS 
 tpg|BK006941.2| 1054486 + tpg|BK006941.2| 1054921 - INS 
 tpg|BK006938.2| 1514710 + tpg|BK006938.2| 1514307 - INS 
 tpg|BK006941.2| 606351 + tpg|BK006941.2| 606543 - INS TGAAC
 tpg|BK006941.2| 695041 + tpg|BK006941.2| 695211 - INS 
 tpg|BK006941.2| 35429 + tpg|BK006941.2| 34923 - INS 
 tpg|BK006938.2| 714540 + tpg|BK006938.2| 714108 - INS 
 tpg|BK006938.2| 928718 + tpg|BK006938.2| 928186 - INS 
 tpg|BK006941.2| 648998 + tpg|BK006941.2| 649016 - INS 
 tpg|BK006938.2| 681487 + tpg|BK006938.2| 681324 - INS 
 tpg|BK006941.2| 437968 + tpg|BK006941.2| 437919 - INS 
 tpg|BK006941.2| 347473 + tpg|BK006941.2| 347185 - INS 
 tpg|BK006938.2| 1168058 + tpg|BK006938.2| 1168687 - INS 
 tpg|BK006941.2| 500526 + tpg|BK006941.2| 499917 - INS 
 tpg|BK006941.2| 581334 + tpg|BK006941.2| 581242 - INS 
 tpg|BK006938.2| 679956 + tpg|BK006938.2| 680459 - INS 
 tpg|BK006941.2| 702647 + tpg|BK006941.2| 702389 - INS 
 tpg|BK006941.2| 772784 + tpg|BK006941.2| 772680 - INS 
 tpg|BK006941.2| 957272 + tpg|BK006941.2| 956544 - INS 
 tpg|BK006941.2| 444240 + tpg|BK006941.2| 443912 - INS 
 tpg|BK006941.2| 148158 + tpg|BK006941.2| 148208 - INS 
 tpg|BK006938.2| 622012 + tpg|BK006938.2| 621407 - INS 
 tpg|BK006941.2| 145511 + tpg|BK006941.2| 145126 - INS 
 tpg|BK006938.2| 245612 + tpg|BK006938.2| 245626 - INS TCAC
 tpg|BK006941.2| 425268 + tpg|BK006941.2| 424804 - INS 
 tpg|BK006938.2| 307771 + tpg|BK006938.2| 307318 - INS 
 tpg|BK006941.2| 797824 + tpg|BK006941.2| 797925 - INS 
 tpg|BK006941.2| 663294 + tpg|BK006941.2| 663920 - INS 
 tpg|BK006941.2| 204855 + tpg|BK006941.2| 204845 - INS 
 tpg|BK006938.2| 915916 + tpg|BK006938.2| 915541 - INS 
 tpg|BK006941.2| 1016428 + tpg|BK006941.2| 1016085 - INS 
 tpg|BK006941.2| 103671 + tpg|BK006941.2| 103631 - INS 
 tpg|BK006938.2| 1001387 + tpg|BK006938.2| 1000667 - INS 
 tpg|BK006941.2| 486497 + tpg|BK006941.2| 486413 - INS 
 tpg|BK006941.2| 969601 + tpg|BK006941.2| 969556 - INS 
 tpg|BK006941.2| 706708 + tpg|BK006941.2| 706273 - INS 
 tpg|BK006941.2| 439224 + tpg|BK006941.2| 439710 - INS 
 tpg|BK006941.2| 318860 + tpg|BK006941.2| 319627 - INS 
 tpg|BK006941.2| 698424 + tpg|BK006941.2| 698720 - INS 
 tpg|BK006941.2| 233638 + tpg|BK006941.2| 233249 - INS 
 tpg|BK006941.2| 685635 + tpg|BK006941.2| 685292 - INS 
 tpg|BK006941.2| 131626 + tpg|BK006941.2| 131928 - INS 
 tpg|BK006941.2| 834848 + tpg|BK006941.2| 834849 - INS 
 tpg|BK006941.2| 37913 + tpg|BK006941.2| 37869 - INS 
 tpg|BK006941.2| 178274 + tpg|BK006941.2| 178131 - INS 
 tpg|BK006941.2| 989695 + tpg|BK006941.2| 989658 - INS 
 tpg|BK006938.2| 1464301 + tpg|BK006938.2| 1463778 - INS 
 tpg|BK006938.2| 190900 + tpg|BK006938.2| 190244 - INS 
 tpg|BK006941.2| 1029165 + tpg|BK006941.2| 1028567 - INS 
 tpg|BK006941.2| 466263 + tpg|BK006941.2| 465823 - INS 
 tpg|BK006941.2| 176491 + tpg|BK006941.2| 176883 - INS 
 tpg|BK006938.2| 300991 + tpg|BK006938.2| 300599 - INS 
 tpg|BK006941.2| 708447 + tpg|BK006941.2| 708155 - INS 
 tpg|BK006941.2| 798941 + tpg|BK006941.2| 798574 - INS 
 tpg|BK006941.2| 686968 + tpg|BK006941.2| 686560 - INS 
 tpg|BK006938.2| 1433797 + tpg|BK006938.2| 1433437 - INS 
 tpg|BK006941.2| 805919 + tpg|BK006941.2| 805489 - INS 
 tpg|BK006941.2| 535747 + tpg|BK006941.2| 535472 - INS 
 tpg|BK006938.2| 1426317 + tpg|BK006938.2| 1425819 - INS 
 tpg|BK006941.2| 791552 + tpg|BK006941.2| 792252 - INS 
 tpg|BK006941.2| 497195 + tpg|BK006941.2| 496879 - INS 
 tpg|BK006941.2| 490866 + tpg|BK006941.2| 491166 - INS 
 tpg|BK006938.2| 266004 + tpg|BK006938.2| 265886 - INS 
 tpg|BK006941.2| 712931 + tpg|BK006941.2| 712474 - INS 
 tpg|BK006941.2| 899867 + tpg|BK006941.2| 899449 - INS 
 tpg|BK006938.2| 585839 + tpg|BK006938.2| 585940 - INS 
 tpg|BK006941.2| 46797 + tpg|BK006941.2| 46200 - INS 
 tpg|BK006941.2| 487389 + tpg|BK006941.2| 486852 - INS 
 tpg|BK006941.2| 222622 + tpg|BK006941.2| 223127 - INS 
 tpg|BK006941.2| 688065 + tpg|BK006941.2| 687560 - INS 
 tpg|BK006941.2| 919113 + tpg|BK006941.2| 919576 - INS 
 tpg|BK006938.2| 148530 + tpg|BK006938.2| 148448 - INS 
 tpg|BK006941.2| 181906 + tpg|BK006941.2| 181735 - INS 
 tpg|BK006941.2| 913073 + tpg|BK006941.2| 912794 - INS 
 tpg|BK006941.2| 216595 + tpg|BK006941.2| 216561 - INS 
 tpg|BK006938.2| 1056641 + tpg|BK006938.2| 1056305 - INS 
 tpg|BK006941.2| 403577 + tpg|BK006941.2| 403311 - INS 
 tpg|BK006938.2| 1066672 + tpg|BK006938.2| 1066268 - INS 
 tpg|BK006938.2| 1109537 + tpg|BK006938.2| 1109143 - INS 
 tpg|BK006938.2| 492459 + tpg|BK006938.2| 491965 - INS 
 tpg|BK006938.2| 1177858 + tpg|BK006938.2| 1178508 - INS 
 tpg|BK006938.2| 1223452 + tpg|BK006938.2| 1223278 - INS 
 tpg|BK006938.2| 321054 + tpg|BK006938.2| 321681 - INS 
 tpg|BK006938.2| 175038 + tpg|BK006938.2| 175028 - INS 
 tpg|BK006938.2| 1372860 + tpg|BK006938.2| 1372782 - INS 
 tpg|BK006938.2| 329016 + tpg|BK006938.2| 328851 - INS 
 tpg|BK006938.2| 1281248 + tpg|BK006938.2| 1281038 - INS 
 tpg|BK006938.2| 1288136 + tpg|BK006938.2| 1288357 - INS 
 tpg|BK006938.2| 336984 + tpg|BK006938.2| 337195 - INS 
 tpg|BK006938.2| 350953 + tpg|BK006938.2| 351025 - INS 
 tpg|BK006938.2| 1335195 + tpg|BK006938.2| 1335892 - INS 
 tpg|BK006938.2| 1145048 + tpg|BK006938.2| 1144301 - INS 
 tpg|BK006938.2| 773491 + tpg|BK006938.2| 773417 - INS 
 tpg|BK006938.2| 808033 + tpg|BK006938.2| 807394 - INS 
 tpg|BK006938.2| 1509688 + tpg|BK006938.2| 1510015 - INS 
 tpg|BK006938.2| 796718 + tpg|BK006938.2| 796170 - INS 
 tpg|BK006938.2| 1508714 + tpg|BK006938.2| 1508089 - INS 
 tpg|BK006938.2| 1469983 + tpg|BK006938.2| 1469843 - INS 
 tpg|BK006938.2| 981299 + tpg|BK006938.2| 980579 - INS 
 tpg|BK006938.2| 372057 + tpg|BK006938.2| 372766 - INS 
 tpg|BK006938.2| 810562 + tpg|BK006938.2| 810648 - INS 
 tpg|BK006938.2| 392071 + tpg|BK006938.2| 392110 - INS 
 tpg|BK006938.2| 631041 + tpg|BK006938.2| 630676 - INS 
 tpg|BK006938.2| 630595 + tpg|BK006938.2| 629945 - INS 
 tpg|BK006938.2| 1090807 + tpg|BK006938.2| 1090195 - INS 
 tpg|BK006938.2| 137231 + tpg|BK006938.2| 137389 - INS 
 tpg|BK006938.2| 581220 + tpg|BK006938.2| 581962 - INS 
 tpg|BK006938.2| 1108462 + tpg|BK006938.2| 1108635 - INS 
 tpg|BK006938.2| 578307 + tpg|BK006938.2| 578017 - INS 
 tpg|BK006938.2| 1305062 + tpg|BK006938.2| 1305768 - INS 
 tpg|BK006938.2| 573913 + tpg|BK006938.2| 574675 - INS 
 tpg|BK006938.2| 890257 + tpg|BK006938.2| 889544 - INS 
 tpg|BK006938.2| 1132827 + tpg|BK006938.2| 1132304 - INS 
 tpg|BK006938.2| 89610 + tpg|BK006938.2| 90102 - INS 
 tpg|BK006938.2| 925522 + tpg|BK006938.2| 925373 - INS 
 tpg|BK006938.2| 619219 + tpg|BK006938.2| 618564 - INS 
 tpg|BK006938.2| 964829 + tpg|BK006938.2| 964803 - INS 
 tpg|BK006938.2| 1393222 + tpg|BK006938.2| 1392882 - INS 
 tpg|BK006938.2| 635508 + tpg|BK006938.2| 635050 - INS 
 tpg|BK006938.2| 452469 + tpg|BK006938.2| 452584 - INS 
 tpg|BK006938.2| 444901 + tpg|BK006938.2| 445224 - INS 
 tpg|BK006938.2| 1153697 + tpg|BK006938.2| 1153654 - INS 
 tpg|BK006938.2| 1444167 + tpg|BK006938.2| 1444806 - INS 
 tpg|BK006938.2| 388429 + tpg|BK006938.2| 388291 - INS 
 tpg|BK006938.2| 687054 + tpg|BK006938.2| 686675 - INS 
 tpg|BK006938.2| 418860 + tpg|BK006938.2| 419165 - INS 
 tpg|BK006938.2| 1152366 + tpg|BK006938.2| 1152263 - INS 
 tpg|BK006938.2| 393031 + tpg|BK006938.2| 392854 - INS 
 tpg|BK006938.2| 389814 + tpg|BK006938.2| 389341 - INS 
 tpg|BK006938.2| 54907 + tpg|BK006938.2| 55160 - INS 
 tpg|BK006938.2| 917973 + tpg|BK006938.2| 918257 - INS 
 tpg|BK006938.2| 197343 + tpg|BK006938.2| 197005 - INS 
 tpg|BK006938.2| 383242 + tpg|BK006938.2| 383381 - INS 
 tpg|BK006938.2| 1250689 + tpg|BK006938.2| 1250511 - INS 
 tpg|BK006938.2| 828356 + tpg|BK006938.2| 827919 - INS 
 tpg|BK006938.2| 742046 + tpg|BK006938.2| 742609 - INS 
 tpg|BK006938.2| 1480717 + tpg|BK006938.2| 1480556 - INS 
 tpg|BK006938.2| 672284 + tpg|BK006938.2| 672838 - INS 
 tpg|BK006938.2| 431178 + tpg|BK006938.2| 431396 - INS 
 tpg|BK006938.2| 918681 + tpg|BK006938.2| 919106 - INS 
 tpg|BK006938.2| 1198710 + tpg|BK006938.2| 1198864 - INS 
 tpg|BK006938.2| 172904 + tpg|BK006938.2| 173513 - INS 
 tpg|BK006938.2| 248459 + tpg|BK006938.2| 248017 - INS 
 tpg|BK006938.2| 660498 + tpg|BK006938.2| 660608 - INS 
 tpg|BK006938.2| 1391531 + tpg|BK006938.2| 1390794 - INS 
 tpg|BK006938.2| 909346 + tpg|BK006938.2| 910035 - INS 
 tpg|BK006938.2| 736146 + tpg|BK006938.2| 736736 - INS 
 tpg|BK006938.2| 932022 + tpg|BK006938.2| 931587 - INS 
 tpg|BK006938.2| 662841 + tpg|BK006938.2| 662262 - INS 
 tpg|BK006938.2| 453232 + tpg|BK006938.2| 453245 - INS 
 tpg|BK006938.2| 93804 + tpg|BK006938.2| 94318 - INS 
 tpg|BK006938.2| 952556 + tpg|BK006938.2| 952834 - INS 
 tpg|BK006938.2| 459717 + tpg|BK006938.2| 458997 - INS 
 tpg|BK006938.2| 1165451 + tpg|BK006938.2| 1165077 - INS 
 tpg|BK006938.2| 1315705 + tpg|BK006938.2| 1314976 - INS 
 tpg|BK006938.2| 469187 + tpg|BK006938.2| 468470 - INS 
 tpg|BK006938.2| 606842 + tpg|BK006938.2| 607104 - INS 
 tpg|BK006938.2| 1148195 + tpg|BK006938.2| 1147799 - INS 
 tpg|BK006938.2| 495910 + tpg|BK006938.2| 495286 - INS 
 tpg|BK006938.2| 1040348 + tpg|BK006938.2| 1039636 - INS 
 tpg|BK006938.2| 278245 + tpg|BK006938.2| 278181 - INS 
 tpg|BK006938.2| 1125089 + tpg|BK006938.2| 1124535 - INS 
 tpg|BK006938.2| 505393 + tpg|BK006938.2| 505466 - INS 
 tpg|BK006938.2| 1117382 + tpg|BK006938.2| 1117806 - INS 
 tpg|BK006938.2| 567370 + tpg|BK006938.2| 566884 - INS 
 tpg|BK006938.2| 1062018 + tpg|BK006938.2| 1062667 - INS 
 tpg|BK006938.2| 1125871 + tpg|BK006938.2| 1125633 - INS 
 tpg|BK006938.2| 153276 + tpg|BK006938.2| 152788 - INS 
 tpg|BK006938.2| 1490131 + tpg|BK006938.2| 1489550 - INS 
 tpg|BK006938.2| 1438527 + tpg|BK006938.2| 1439077 - INS 
 tpg|BK006938.2| 1394068 + tpg|BK006938.2| 1393450 - INS 
 tpg|BK006938.2| 939397 + tpg|BK006938.2| 939285 - INS 
 tpg|BK006938.2| 1345571 + tpg|BK006938.2| 1344947 - INS 
 tpg|BK006938.2| 467548 + tpg|BK006938.2| 467786 - INS 
 tpg|BK006938.2| 353513 + tpg|BK006938.2| 353283 - INS 
 tpg|BK006938.2| 338131 + tpg|BK006938.2| 338332 - INS 
 tpg|BK006946.2| 759232 + tpg|BK006946.2| 759681 - INS 
 tpg|BK006938.2| 1364111 + tpg|BK006938.2| 1364027 - INS 
 tpg|BK006938.2| 1322767 + tpg|BK006938.2| 1323069 - INS 
 tpg|BK006938.2| 1320173 + tpg|BK006938.2| 1319636 - INS 
 tpg|BK006938.2| 750991 + tpg|BK006938.2| 750482 - INS 
 tpg|BK006946.2| 868810 + tpg|BK006946.2| 869257 - INS 
 tpg|BK006938.2| 1825 + tpg|BK006938.2| 1523 - INS 
 tpg|BK006938.2| 1280530 + tpg|BK006938.2| 1279873 - INS 
 tpg|BK006938.2| 789751 + tpg|BK006938.2| 789444 - INS 
 tpg|BK006938.2| 762999 + tpg|BK006938.2| 762355 - INS 
 tpg|BK006938.2| 809070 + tpg|BK006938.2| 809491 - INS 
 tpg|BK006946.2| 70443 + tpg|BK006946.2| 69857 - INS 
 tpg|BK006938.2| 821887 + tpg|BK006938.2| 821318 - INS 
 tpg|BK006938.2| 741267 + tpg|BK006938.2| 740723 - INS 
 tpg|BK006946.2| 612474 + tpg|BK006946.2| 612587 - INS 
 tpg|BK006938.2| 201416 + tpg|BK006938.2| 202066 - INS 
 tpg|BK006938.2| 1515744 + tpg|BK006938.2| 1515672 - INS 
 tpg|BK006938.2| 676042 + tpg|BK006938.2| 675361 - INS 
 tpg|BK006946.2| 101496 + tpg|BK006946.2| 101972 - INS 
 tpg|BK006938.2| 996765 + tpg|BK006938.2| 997516 - INS 
 tpg|BK006938.2| 1442897 + tpg|BK006938.2| 1442164 - INS 
 tpg|BK006938.2| 1029212 + tpg|BK006938.2| 1029601 - INS 
 tpg|BK006938.2| 587799 + tpg|BK006938.2| 588037 - INS 
 tpg|BK006946.2| 40027 + tpg|BK006946.2| 39374 - INS 
 tpg|BK006938.2| 1052853 + tpg|BK006938.2| 1053601 - INS 
 tpg|BK006938.2| 1067347 + tpg|BK006938.2| 1066868 - INS 
 tpg|BK006946.2| 222765 + tpg|BK006946.2| 222902 - INS 
 tpg|BK006938.2| 1423154 + tpg|BK006938.2| 1423736 - INS 
 tpg|BK006938.2| 1123523 + tpg|BK006938.2| 1122762 - INS 
 tpg|BK006938.2| 1413522 + tpg|BK006938.2| 1413708 - INS 
 tpg|BK006938.2| 29840 + tpg|BK006938.2| 29732 - INS 
 tpg|BK006938.2| 73831 + tpg|BK006938.2| 73387 - INS 
 tpg|BK006938.2| 1032169 + tpg|BK006938.2| 1032294 - INS 
 tpg|BK006946.2| 308288 + tpg|BK006946.2| 308748 - INS 
 tpg|BK006938.2| 507331 + tpg|BK006938.2| 507499 - INS 
 tpg|BK006938.2| 497547 + tpg|BK006938.2| 497361 - INS 
 tpg|BK006938.2| 1398226 + tpg|BK006938.2| 1397500 - INS 
 tpg|BK006946.2| 16716 + tpg|BK006946.2| 16129 - INS 
 tpg|BK006938.2| 1167010 + tpg|BK006938.2| 1166553 - INS 
 tpg|BK006946.2| 660472 + tpg|BK006946.2| 661091 - INS 
 tpg|BK006946.2| 491884 + tpg|BK006946.2| 492180 - INS 
 tpg|BK006946.2| 742763 + tpg|BK006946.2| 742994 - INS 
 tpg|BK006938.2| 966056 + tpg|BK006938.2| 965427 - INS 
 tpg|BK006946.2| 872497 + tpg|BK006946.2| 872356 - INS 
 tpg|BK006938.2| 937709 + tpg|BK006938.2| 937498 - INS 
 tpg|BK006938.2| 1265900 + tpg|BK006938.2| 1266242 - INS 
 tpg|BK006938.2| 1186808 + tpg|BK006938.2| 1187127 - INS 
 tpg|BK006946.2| 334335 + tpg|BK006946.2| 334515 - INS 
 tpg|BK006938.2| 641524 + tpg|BK006938.2| 640987 - INS 
 tpg|BK006938.2| 642971 + tpg|BK006938.2| 642323 - INS 
 tpg|BK006946.2| 41343 + tpg|BK006946.2| 41935 - INS 
 tpg|BK006938.2| 645121 + tpg|BK006938.2| 644413 - INS 
 tpg|BK006938.2| 1285750 + tpg|BK006938.2| 1285274 - INS 
 tpg|BK006946.2| 276509 + tpg|BK006946.2| 275748 - INS 
 tpg|BK006938.2| 430298 + tpg|BK006938.2| 429952 - INS 
 tpg|BK006938.2| 240482 + tpg|BK006938.2| 240106 - INS 
 tpg|BK006938.2| 1353863 + tpg|BK006938.2| 1353707 - INS 
 tpg|BK006938.2| 417943 + tpg|BK006938.2| 418177 - INS 
 tpg|BK006946.2| 763738 + tpg|BK006946.2| 763795 - INS 
 tpg|BK006938.2| 697482 + tpg|BK006938.2| 696775 - INS 
 tpg|BK006938.2| 701717 + tpg|BK006938.2| 701290 - INS 
 tpg|BK006938.2| 231962 + tpg|BK006938.2| 232313 - INS 
 tpg|BK006938.2| 855337 + tpg|BK006938.2| 855406 - INS 
 tpg|BK006946.2| 390356 + tpg|BK006946.2| 389782 - INS 
 tpg|BK006938.2| 393655 + tpg|BK006938.2| 393724 - INS 
 tpg|BK006946.2| 408660 + tpg|BK006946.2| 408578 - INS 
 tpg|BK006938.2| 723346 + tpg|BK006938.2| 722955 - INS 
 tpg|BK006938.2| 735345 + tpg|BK006938.2| 735305 - INS 
 tpg|BK006946.2| 271015 + tpg|BK006946.2| 270935 - INS 
 tpg|BK006938.2| 213169 + tpg|BK006938.2| 213648 - INS 
 tpg|BK006938.2| 1316338 + tpg|BK006938.2| 1315673 - INS 
 tpg|BK006946.2| 316081 + tpg|BK006946.2| 316577 - INS 
 tpg|BK006938.2| 760138 + tpg|BK006938.2| 760721 - INS 
 tpg|BK006938.2| 244394 + tpg|BK006938.2| 244811 - INS 
 tpg|BK006938.2| 998490 + tpg|BK006938.2| 998680 - INS 
 tpg|BK006938.2| 771810 + tpg|BK006938.2| 772249 - INS 
 tpg|BK006946.2| 531043 + tpg|BK006946.2| 530662 - INS 
 tpg|BK006938.2| 1506981 + tpg|BK006938.2| 1506914 - INS 
 tpg|BK006938.2| 1495828 + tpg|BK006938.2| 1495940 - INS 
 tpg|BK006946.2| 884939 + tpg|BK006946.2| 885075 - INS 
 tpg|BK006938.2| 249467 + tpg|BK006938.2| 249796 - INS 
 tpg|BK006938.2| 1436969 + tpg|BK006938.2| 1437133 - INS 
 tpg|BK006938.2| 935875 + tpg|BK006938.2| 936603 - INS 
 tpg|BK006946.2| 367771 + tpg|BK006946.2| 368544 - INS 
 tpg|BK006938.2| 747881 + tpg|BK006938.2| 747947 - INS 
 tpg|BK006946.2| 747560 + tpg|BK006946.2| 747058 - INS 
 tpg|BK006938.2| 397661 + tpg|BK006938.2| 397543 - INS 
 tpg|BK006938.2| 1239253 + tpg|BK006938.2| 1239540 - INS 
 tpg|BK006946.2| 836781 + tpg|BK006946.2| 836694 - INS 
 tpg|BK006946.2| 30379 + tpg|BK006946.2| 29762 - INS 
 tpg|BK006938.2| 812914 + tpg|BK006938.2| 812926 - INS 
 tpg|BK006938.2| 1180904 + tpg|BK006938.2| 1180621 - INS 
 tpg|BK006946.2| 258376 + tpg|BK006946.2| 257714 - INS 
 tpg|BK006946.2| 167121 + tpg|BK006946.2| 166435 - INS 
 tpg|BK006938.2| 891927 + tpg|BK006938.2| 891588 - INS 
 tpg|BK006938.2| 547336 + tpg|BK006938.2| 547352 - INS 
 tpg|BK006946.2| 136883 + tpg|BK006946.2| 137641 - INS 
 tpg|BK006938.2| 926269 + tpg|BK006938.2| 925969 - INS 
 tpg|BK006938.2| 1388842 + tpg|BK006938.2| 1388717 - INS 
 tpg|BK006938.2| 95162 + tpg|BK006938.2| 95015 - INS 
 tpg|BK006938.2| 1231608 + tpg|BK006938.2| 1231287 - INS 
 tpg|BK006938.2| 369576 + tpg|BK006938.2| 369464 - INS 
 tpg|BK006946.2| 659654 + tpg|BK006946.2| 660115 - INS 
 tpg|BK006938.2| 274888 + tpg|BK006938.2| 274161 - INS 
 tpg|BK006938.2| 271493 + tpg|BK006938.2| 271340 - INS 
 tpg|BK006946.2| 657040 + tpg|BK006946.2| 656373 - INS 
 tpg|BK006938.2| 1346375 + tpg|BK006938.2| 1345773 - INS 
 tpg|BK006946.2| 900334 + tpg|BK006946.2| 900992 - INS 
 tpg|BK006946.2| 220807 + tpg|BK006946.2| 220324 - INS 
 tpg|BK006938.2| 1263598 + tpg|BK006938.2| 1264278 - INS 
 tpg|BK006938.2| 863575 + tpg|BK006938.2| 863585 - INS 
 tpg|BK006938.2| 1257364 + tpg|BK006938.2| 1257714 - INS 
 tpg|BK006938.2| 885283 + tpg|BK006938.2| 884750 - INS 
 tpg|BK006938.2| 65728 + tpg|BK006938.2| 65264 - INS 
 tpg|BK006946.2| 473970 + tpg|BK006946.2| 474671 - INS 
 tpg|BK006938.2| 434465 + tpg|BK006938.2| 434953 - INS 
 tpg|BK006938.2| 639945 + tpg|BK006938.2| 639408 - INS 
 tpg|BK006938.2| 1461481 + tpg|BK006938.2| 1461307 - INS 
 tpg|BK006938.2| 1182477 + tpg|BK006938.2| 1181712 - INS 
 tpg|BK006946.2| 278317 + tpg|BK006946.2| 278124 - INS 
 tpg|BK006938.2| 1179422 + tpg|BK006938.2| 1179117 - INS 
 tpg|BK006938.2| 1174975 + tpg|BK006938.2| 1174648 - INS 
 tpg|BK006946.2| 445278 + tpg|BK006946.2| 444945 - INS 
 tpg|BK006938.2| 165894 + tpg|BK006938.2| 166500 - INS 
 tpg|BK006938.2| 93240 + tpg|BK006938.2| 93042 - INS 
 tpg|BK006946.2| 219008 + tpg|BK006946.2| 219710 - INS 
 tpg|BK006938.2| 1185523 + tpg|BK006938.2| 1185288 - INS 
 tpg|BK006946.2| 673934 + tpg|BK006946.2| 673883 - INS 
 tpg|BK006938.2| 616286 + tpg|BK006938.2| 615949 - INS 
 tpg|BK006938.2| 1163086 + tpg|BK006938.2| 1162690 - INS 
 tpg|BK006938.2| 263353 + tpg|BK006938.2| 262773 - INS 
 tpg|BK006946.2| 820556 + tpg|BK006946.2| 820249 - INS 
 tpg|BK006938.2| 546603 + tpg|BK006938.2| 545882 - INS 
 tpg|BK006946.2| 479273 + tpg|BK006946.2| 479412 - INS 
 tpg|BK006938.2| 1443389 + tpg|BK006938.2| 1443283 - INS 
 tpg|BK006946.2| 363306 + tpg|BK006946.2| 363344 - INS 
 tpg|BK006946.2| 110363 + tpg|BK006946.2| 110531 - INS 
 tpg|BK006938.2| 83580 + tpg|BK006938.2| 84347 - INS 
 tpg|BK006938.2| 1149181 + tpg|BK006938.2| 1148537 - INS 
 tpg|BK006938.2| 1048954 + tpg|BK006938.2| 1048552 - INS 
 tpg|BK006946.2| 797479 + tpg|BK006946.2| 797397 - INS 
 tpg|BK006938.2| 31315 + tpg|BK006938.2| 31535 - INS 
 tpg|BK006938.2| 186036 + tpg|BK006938.2| 186487 - INS 
 tpg|BK006938.2| 1064741 + tpg|BK006938.2| 1064718 - INS 
 tpg|BK006946.2| 875250 + tpg|BK006946.2| 875098 - INS 
 tpg|BK006938.2| 1111627 + tpg|BK006938.2| 1111157 - INS 
 tpg|BK006946.2| 560052 + tpg|BK006946.2| 560723 - INS 
 tpg|BK006938.2| 541342 + tpg|BK006938.2| 541075 - INS 
 tpg|BK006938.2| 552795 + tpg|BK006938.2| 552739 - INS 
 tpg|BK006938.2| 1412634 + tpg|BK006938.2| 1412216 - INS 
 tpg|BK006938.2| 1092659 + tpg|BK006938.2| 1093341 - INS 
 tpg|BK006938.2| 1350132 + tpg|BK006938.2| 1350724 - INS 
 tpg|BK006938.2| 1118773 + tpg|BK006938.2| 1119168 - INS 
 tpg|BK006938.2| 1426907 + tpg|BK006938.2| 1426764 - INS 
 tpg|BK006946.2| 808506 + tpg|BK006946.2| 808282 - INS 
 tpg|BK006938.2| 1031358 + tpg|BK006938.2| 1030831 - INS 
 tpg|BK006938.2| 1402766 + tpg|BK006938.2| 1402738 - INS 
 tpg|BK006946.2| 344992 + tpg|BK006946.2| 344855 - INS 
 tpg|BK006938.2| 590469 + tpg|BK006938.2| 590127 - INS 
 tpg|BK006938.2| 1029610 + tpg|BK006938.2| 1030279 - INS 
 tpg|BK006946.2| 209083 + tpg|BK006946.2| 209148 - INS 
 tpg|BK006938.2| 591355 + tpg|BK006938.2| 591209 - INS 
 tpg|BK006946.2| 170810 + tpg|BK006946.2| 170045 - INS 
 tpg|BK006938.2| 305967 + tpg|BK006938.2| 305919 - INS 
 tpg|BK006938.2| 1008945 + tpg|BK006938.2| 1009465 - INS 
 tpg|BK006946.2| 754885 + tpg|BK006946.2| 754299 - INS 
 tpg|BK006946.2| 135125 + tpg|BK006946.2| 135090 - INS 
 tpg|BK006938.2| 470162 + tpg|BK006938.2| 469797 - INS 
 tpg|BK006938.2| 969259 + tpg|BK006938.2| 968883 - INS 
 tpg|BK006946.2| 715131 + tpg|BK006946.2| 715068 - INS 
 tpg|BK006946.2| 768255 + tpg|BK006946.2| 767858 - INS 
 tpg|BK006946.2| 623662 + tpg|BK006946.2| 622991 - INS 
 tpg|BK006938.2| 963897 + tpg|BK006938.2| 963755 - INS 
 tpg|BK006938.2| 1166303 + tpg|BK006938.2| 1165952 - INS 
 tpg|BK006938.2| 628921 + tpg|BK006938.2| 628483 - INS 
 tpg|BK006946.2| 778751 + tpg|BK006946.2| 778143 - INS 
 tpg|BK006946.2| 280741 + tpg|BK006946.2| 280687 - INS 
 tpg|BK006938.2| 441211 + tpg|BK006938.2| 441241 - INS 
 tpg|BK006938.2| 920590 + tpg|BK006938.2| 919861 - INS 
 tpg|BK006938.2| 668651 + tpg|BK006938.2| 669355 - INS 
 tpg|BK006946.2| 451177 + tpg|BK006946.2| 451126 - INS 
 tpg|BK006938.2| 914852 + tpg|BK006938.2| 914742 - INS 
 tpg|BK006938.2| 913638 + tpg|BK006938.2| 913702 - INS 
 tpg|BK006946.2| 272752 + tpg|BK006946.2| 272366 - INS 
 tpg|BK006938.2| 1214833 + tpg|BK006938.2| 1214356 - INS 
 tpg|BK006946.2| 31536 + tpg|BK006946.2| 31075 - INS 
 tpg|BK006938.2| 908301 + tpg|BK006938.2| 907930 - INS 
 tpg|BK006938.2| 673818 + tpg|BK006938.2| 673366 - INS 
 tpg|BK006946.2| 793405 + tpg|BK006946.2| 793399 - INS 
 tpg|BK006938.2| 779553 + tpg|BK006938.2| 779256 - INS 
 tpg|BK006946.2| 608771 + tpg|BK006946.2| 608207 - INS 
 tpg|BK006938.2| 693470 + tpg|BK006938.2| 694116 - INS 
 tpg|BK006946.2| 694591 + tpg|BK006946.2| 694607 - INS 
 tpg|BK006938.2| 777582 + tpg|BK006938.2| 777422 - INS 
 tpg|BK006938.2| 414995 + tpg|BK006938.2| 414707 - INS 
 tpg|BK006938.2| 704023 + tpg|BK006938.2| 704268 - INS 
 tpg|BK006946.2| 372011 + tpg|BK006946.2| 372208 - INS 
 tpg|BK006938.2| 42418 + tpg|BK006938.2| 42348 - INS 
 tpg|BK006938.2| 1256874 + tpg|BK006938.2| 1257046 - INS 
 tpg|BK006938.2| 325192 + tpg|BK006938.2| 325090 - INS 
 tpg|BK006938.2| 220509 + tpg|BK006938.2| 219969 - INS 
 tpg|BK006946.2| 61731 + tpg|BK006946.2| 61386 - INS 
 tpg|BK006938.2| 1300698 + tpg|BK006938.2| 1300801 - INS 
 tpg|BK006938.2| 331321 + tpg|BK006938.2| 331806 - INS 
 tpg|BK006946.2| 124164 + tpg|BK006946.2| 124721 - INS 
 tpg|BK006938.2| 816370 + tpg|BK006938.2| 816629 - INS 
 tpg|BK006938.2| 826303 + tpg|BK006938.2| 826857 - INS 
 tpg|BK006946.2| 860489 + tpg|BK006946.2| 860420 - INS 
 tpg|BK006938.2| 799287 + tpg|BK006938.2| 798670 - INS 
 tpg|BK006938.2| 792219 + tpg|BK006938.2| 791982 - INS 
 tpg|BK006946.2| 454121 + tpg|BK006946.2| 454473 - INS 
 tpg|BK006938.2| 235944 + tpg|BK006938.2| 236101 - INS 
 tpg|BK006946.2| 447656 + tpg|BK006946.2| 447968 - INS 
 tpg|BK006938.2| 794648 + tpg|BK006938.2| 793905 - INS 
 tpg|BK006938.2| 758047 + tpg|BK006938.2| 757274 - INS 
 tpg|BK006946.2| 250238 + tpg|BK006946.2| 250239 - INS 
 tpg|BK006938.2| 832331 + tpg|BK006938.2| 831839 - INS 
 tpg|BK006938.2| 222965 + tpg|BK006938.2| 223298 - INS 
 tpg|BK006938.2| 1406608 + tpg|BK006938.2| 1406906 - INS 
 tpg|BK006946.2| 12488 + tpg|BK006946.2| 11980 - INS 
 tpg|BK006938.2| 301692 + tpg|BK006938.2| 301274 - INS 
 tpg|BK006946.2| 662564 + tpg|BK006946.2| 662833 - INS 
 tpg|BK006938.2| 34573 + tpg|BK006938.2| 34865 - INS 
 tpg|BK006938.2| 869286 + tpg|BK006938.2| 869839 - INS 
 tpg|BK006946.2| 583970 + tpg|BK006946.2| 583832 - INS 
 tpg|BK006938.2| 670060 + tpg|BK006938.2| 670004 - INS 
 tpg|BK006946.2| 65316 + tpg|BK006946.2| 65851 - INS 
 tpg|BK006938.2| 1360063 + tpg|BK006938.2| 1359602 - INS 
 tpg|BK006946.2| 205947 + tpg|BK006946.2| 206234 - INS 
 tpg|BK006938.2| 922968 + tpg|BK006938.2| 922453 - INS 
 tpg|BK006946.2| 515298 + tpg|BK006946.2| 516040 - INS 
 tpg|BK006938.2| 1494937 + tpg|BK006938.2| 1494939 - INS 
 tpg|BK006946.2| 326680 + tpg|BK006946.2| 326364 - INS 
 tpg|BK006938.2| 1493565 + tpg|BK006938.2| 1493084 - INS 
 tpg|BK006946.2| 468274 + tpg|BK006946.2| 468272 - INS 
 tpg|BK006938.2| 1309058 + tpg|BK006938.2| 1308527 - INS 
 tpg|BK006938.2| 251383 + tpg|BK006938.2| 251378 - INS 
 tpg|BK006946.2| 338028 + tpg|BK006946.2| 337761 - INS 
 tpg|BK006938.2| 133776 + tpg|BK006938.2| 134042 - INS 
 tpg|BK006938.2| 1467486 + tpg|BK006938.2| 1467099 - INS 
 tpg|BK006938.2| 409709 + tpg|BK006938.2| 409299 - INS 
 tpg|BK006938.2| 1008231 + tpg|BK006938.2| 1007967 - INS 
 tpg|BK006938.2| 1012240 + tpg|BK006938.2| 1012990 - INS 
 tpg|BK006938.2| 447188 + tpg|BK006938.2| 446920 - INS 
 tpg|BK006938.2| 975411 + tpg|BK006938.2| 975103 - INS 
 tpg|BK006938.2| 611457 + tpg|BK006938.2| 610743 - INS 
 tpg|BK006946.2| 745249 + tpg|BK006946.2| 745043 - INS 
 tpg|BK006946.2| 405411 + tpg|BK006946.2| 405341 - INS 
 tpg|BK006938.2| 998995 + tpg|BK006938.2| 999276 - INS 
 tpg|BK006946.2| 710069 + tpg|BK006946.2| 710259 - INS 
 tpg|BK006938.2| 82606 + tpg|BK006938.2| 82757 - INS 
 tpg|BK006946.2| 716339 + tpg|BK006946.2| 716130 - INS 
 tpg|BK006938.2| 540466 + tpg|BK006938.2| 539711 - INS 
 tpg|BK006946.2| 406993 + tpg|BK006946.2| 407242 - INS 
 tpg|BK006938.2| 1110645 + tpg|BK006938.2| 1110370 - INS 
 tpg|BK006938.2| 1046652 + tpg|BK006938.2| 1046280 - INS 
 tpg|BK006946.2| 402072 + tpg|BK006946.2| 401748 - INS 
 tpg|BK006938.2| 1047430 + tpg|BK006938.2| 1046756 - INS 
 tpg|BK006938.2| 1084330 + tpg|BK006938.2| 1083871 - INS 
 tpg|BK006938.2| 503583 + tpg|BK006938.2| 503087 - INS 
 tpg|BK006938.2| 171549 + tpg|BK006938.2| 171281 - INS 
 tpg|BK006938.2| 1271211 + tpg|BK006938.2| 1270876 - INS 
 tpg|BK006946.2| 178485 + tpg|BK006946.2| 178641 - INS 
 tpg|BK006938.2| 1295127 + tpg|BK006938.2| 1295053 - INS 
 tpg|BK006938.2| 183417 + tpg|BK006938.2| 183269 - INS 
 tpg|BK006938.2| 852355 + tpg|BK006938.2| 852638 - INS 
 tpg|BK006946.2| 14250 + tpg|BK006946.2| 14415 - INS 
 tpg|BK006938.2| 1474219 + tpg|BK006938.2| 1474070 - INS 
 tpg|BK006938.2| 451668 + tpg|BK006938.2| 451633 - INS 
 tpg|BK006946.2| 35124 + tpg|BK006946.2| 35333 - INS 
 tpg|BK006938.2| 429454 + tpg|BK006938.2| 429204 - INS 
 tpg|BK006938.2| 1401400 + tpg|BK006938.2| 1401901 - INS 
 tpg|BK006938.2| 1389996 + tpg|BK006938.2| 1389459 - INS 
 tpg|BK006938.2| 1366529 + tpg|BK006938.2| 1366376 - INS 
 tpg|BK006938.2| 733393 + tpg|BK006938.2| 733529 - INS 
 tpg|BK006938.2| 1086381 + tpg|BK006938.2| 1086933 - INS 
 tpg|BK006938.2| 551832 + tpg|BK006938.2| 552042 - INS 
 tpg|BK006938.2| 1074168 + tpg|BK006938.2| 1073799 - INS 
 tpg|BK006938.2| 1089538 + tpg|BK006938.2| 1089650 - INS 
 tpg|BK006946.2| 658070 + tpg|BK006946.2| 657550 - INS 
 tpg|BK006946.2| 37286 + tpg|BK006946.2| 37587 - INS 
 tpg|BK006938.2| 1050132 + tpg|BK006938.2| 1050168 - INS 
 tpg|BK006946.2| 386735 + tpg|BK006946.2| 386958 - INS 
 tpg|BK006938.2| 146186 + tpg|BK006938.2| 146795 - INS 
 tpg|BK006938.2| 1040944 + tpg|BK006938.2| 1040305 - INS 
 tpg|BK006946.2| 255749 + tpg|BK006946.2| 255159 - INS 
 tpg|BK006938.2| 304496 + tpg|BK006938.2| 305220 - INS 
 tpg|BK006938.2| 1140432 + tpg|BK006938.2| 1139762 - INS 
 tpg|BK006938.2| 70728 + tpg|BK006938.2| 70847 - INS 
 tpg|BK006946.2| 44792 + tpg|BK006946.2| 44514 - INS 
 tpg|BK006938.2| 142957 + tpg|BK006938.2| 142739 - INS 
 tpg|BK006946.2| 172833 + tpg|BK006946.2| 172252 - INS 
 tpg|BK006946.2| 312861 + tpg|BK006946.2| 312512 - INS 
 tpg|BK006938.2| 470862 + tpg|BK006938.2| 470464 - INS 
 tpg|BK006938.2| 994780 + tpg|BK006938.2| 994026 - INS 
 tpg|BK006946.2| 700783 + tpg|BK006946.2| 700528 - INS 
 tpg|BK006938.2| 1453962 + tpg|BK006938.2| 1453343 - INS 
 tpg|BK006938.2| 629734 + tpg|BK006938.2| 629100 - INS 
 tpg|BK006946.2| 817334 + tpg|BK006946.2| 817955 - INS 
 tpg|BK006938.2| 450016 + tpg|BK006938.2| 449356 - INS 
 tpg|BK006938.2| 1466442 + tpg|BK006938.2| 1465705 - INS 
 tpg|BK006946.2| 147684 + tpg|BK006946.2| 147467 - INS 
 tpg|BK006938.2| 1472265 + tpg|BK006938.2| 1472795 - INS 
 tpg|BK006946.2| 45489 + tpg|BK006946.2| 45858 - INS 
 tpg|BK006938.2| 891354 + tpg|BK006938.2| 890889 - INS 
 tpg|BK006938.2| 1230761 + tpg|BK006938.2| 1230086 - INS 
 tpg|BK006946.2| 634155 + tpg|BK006946.2| 633488 - INS 
 tpg|BK006938.2| 1515345 + tpg|BK006938.2| 1514830 - INS 
 tpg|BK006938.2| 854003 + tpg|BK006938.2| 853276 - INS 
 tpg|BK006946.2| 407576 + tpg|BK006946.2| 407878 - INS 
 tpg|BK006938.2| 1270266 + tpg|BK006938.2| 1270063 - INS 
 tpg|BK006946.2| 98901 + tpg|BK006946.2| 98593 - INS 
 tpg|BK006938.2| 729330 + tpg|BK006938.2| 728999 - INS 
 tpg|BK006938.2| 838117 + tpg|BK006938.2| 837710 - INS 
 tpg|BK006946.2| 100878 + tpg|BK006946.2| 100316 - INS 
 tpg|BK006938.2| 330599 + tpg|BK006938.2| 330105 - INS 
 tpg|BK006946.2| 273898 + tpg|BK006946.2| 274645 - INS 
 tpg|BK006946.2| 182036 + tpg|BK006946.2| 181409 - INS 
 tpg|BK006938.2| 1287080 + tpg|BK006938.2| 1287595 - INS 
 tpg|BK006946.2| 248136 + tpg|BK006946.2| 247929 - INS 
 tpg|BK006938.2| 334731 + tpg|BK006938.2| 334118 - INS 
 tpg|BK006938.2| 115718 + tpg|BK006938.2| 115948 - INS 
 tpg|BK006946.2| 750946 + tpg|BK006946.2| 750466 - INS 
 tpg|BK006938.2| 767190 + tpg|BK006938.2| 767533 - INS 
 tpg|BK006938.2| 351932 + tpg|BK006938.2| 351533 - INS 
 tpg|BK006946.2| 548970 + tpg|BK006946.2| 548842 - INS 
 tpg|BK006938.2| 122303 + tpg|BK006938.2| 121639 - INS 
 tpg|BK006938.2| 716890 + tpg|BK006938.2| 716830 - INS 
 tpg|BK006938.2| 716237 + tpg|BK006938.2| 715974 - INS 
 tpg|BK006938.2| 1265234 + tpg|BK006938.2| 1264779 - INS 
 tpg|BK006946.2| 762994 + tpg|BK006946.2| 763054 - INS 
 tpg|BK006938.2| 399777 + tpg|BK006938.2| 399904 - INS 
 tpg|BK006938.2| 400981 + tpg|BK006938.2| 400523 - INS 
 tpg|BK006946.2| 347828 + tpg|BK006946.2| 348562 - INS 
 tpg|BK006938.2| 1262633 + tpg|BK006938.2| 1262165 - INS 
 tpg|BK006938.2| 1259606 + tpg|BK006938.2| 1259906 - INS 
 tpg|BK006946.2| 883439 + tpg|BK006946.2| 883147 - INS 
 tpg|BK006938.2| 1471301 + tpg|BK006938.2| 1470626 - INS 
 tpg|BK006938.2| 1468220 + tpg|BK006938.2| 1468629 - INS 
 tpg|BK006938.2| 1512083 + tpg|BK006938.2| 1511860 - INS 
 tpg|BK006938.2| 254424 + tpg|BK006938.2| 253836 - INS 
 tpg|BK006946.2| 679977 + tpg|BK006946.2| 679540 - INS 
 tpg|BK006938.2| 1458301 + tpg|BK006938.2| 1458326 - INS 
 tpg|BK006938.2| 192547 + tpg|BK006938.2| 192023 - INS 
 tpg|BK006946.2| 324857 + tpg|BK006946.2| 324694 - INS 
 tpg|BK006938.2| 1439467 + tpg|BK006938.2| 1439534 - INS 
 tpg|BK006938.2| 198105 + tpg|BK006938.2| 197883 - INS 
 tpg|BK006946.2| 394607 + tpg|BK006946.2| 394061 - INS 
 tpg|BK006938.2| 1218993 + tpg|BK006938.2| 1219394 - INS 
 tpg|BK006946.2| 410704 + tpg|BK006946.2| 411403 - INS 
 tpg|BK006938.2| 1417434 + tpg|BK006938.2| 1417202 - INS 
 tpg|BK006946.2| 724197 + tpg|BK006946.2| 724916 - INS 
 tpg|BK006938.2| 297983 + tpg|BK006938.2| 297921 - INS 
 tpg|BK006938.2| 894750 + tpg|BK006938.2| 895018 - INS 
 tpg|BK006938.2| 21288 + tpg|BK006938.2| 20997 - INS 
 tpg|BK006938.2| 1370993 + tpg|BK006938.2| 1370330 - INS 
 tpg|BK006946.2| 10697 + tpg|BK006946.2| 10485 - INS 
 tpg|BK006938.2| 1184130 + tpg|BK006938.2| 1183914 - INS 
 tpg|BK006938.2| 1451163 + tpg|BK006938.2| 1451127 - INS 
 tpg|BK006946.2| 346601 + tpg|BK006946.2| 346852 - INS 
 tpg|BK006938.2| 631883 + tpg|BK006938.2| 631871 - INS 
 tpg|BK006938.2| 724410 + tpg|BK006938.2| 725121 - INS 
 tpg|BK006938.2| 1339730 + tpg|BK006938.2| 1339442 - INS 
 tpg|BK006938.2| 193448 + tpg|BK006938.2| 194025 - INS 
 tpg|BK006938.2| 310871 + tpg|BK006938.2| 310454 - INS 
 tpg|BK006946.2| 53707 + tpg|BK006946.2| 53332 - INS 
 tpg|BK006946.2| 141428 + tpg|BK006946.2| 140813 - INS 
 tpg|BK006946.2| 594038 + tpg|BK006946.2| 593366 - INS 
 tpg|BK006938.2| 1362162 + tpg|BK006938.2| 1362296 - INS 
 tpg|BK006946.2| 504553 + tpg|BK006946.2| 504155 - INS 
 tpg|BK006938.2| 136476 + tpg|BK006938.2| 136125 - INS 
 tpg|BK006946.2| 25861 + tpg|BK006946.2| 25779 - INS 
 tpg|BK006938.2| 1298253 + tpg|BK006938.2| 1297517 - INS 
 tpg|BK006938.2| 922161 + tpg|BK006938.2| 921707 - INS 
 tpg|BK006938.2| 549237 + tpg|BK006938.2| 548853 - INS 
 tpg|BK006946.2| 226140 + tpg|BK006946.2| 225368 - INS 
 tpg|BK006938.2| 390333 + tpg|BK006938.2| 390249 - INS GTTATCGTTAT
 tpg|BK006938.2| 1238507 + tpg|BK006938.2| 1238014 - INS 
 tpg|BK006938.2| 416315 + tpg|BK006938.2| 415829 - INS 
 tpg|BK006946.2| 614078 + tpg|BK006946.2| 614004 - INS 
 tpg|BK006938.2| 493612 + tpg|BK006938.2| 493174 - INS 
 tpg|BK006938.2| 1435899 + tpg|BK006938.2| 1435969 - INS 
 tpg|BK006938.2| 1204034 + tpg|BK006938.2| 1203699 - INS 
 tpg|BK006946.2| 723621 + tpg|BK006946.2| 723157 - INS 
 tpg|BK006938.2| 68667 + tpg|BK006938.2| 67958 - INS 
 tpg|BK006946.2| 615955 + tpg|BK006946.2| 616373 - INS 
 tpg|BK006938.2| 1091867 + tpg|BK006938.2| 1091151 - INS 
 tpg|BK006938.2| 521181 + tpg|BK006938.2| 521382 - INS 
 tpg|BK006938.2| 1104848 + tpg|BK006938.2| 1105166 - INS 
 tpg|BK006946.2| 850944 + tpg|BK006946.2| 850382 - INS 
 tpg|BK006938.2| 80518 + tpg|BK006938.2| 80986 - INS 
 tpg|BK006938.2| 204595 + tpg|BK006938.2| 203951 - INS 
 tpg|BK006938.2| 489627 + tpg|BK006938.2| 489823 - INS 
 tpg|BK006938.2| 1070328 + tpg|BK006938.2| 1070207 - INS 
 tpg|BK006946.2| 418048 + tpg|BK006946.2| 418393 - INS 
 tpg|BK006938.2| 153675 + tpg|BK006938.2| 153545 - INS 
 tpg|BK006938.2| 78273 + tpg|BK006938.2| 78291 - INS 
 tpg|BK006946.2| 269889 + tpg|BK006946.2| 270390 - INS 
 tpg|BK006938.2| 1123854 + tpg|BK006938.2| 1123704 - INS 
 tpg|BK006946.2| 104997 + tpg|BK006946.2| 104673 - INS 
 tpg|BK006938.2| 512212 + tpg|BK006938.2| 511734 - INS 
 tpg|BK006946.2| 387376 + tpg|BK006946.2| 387876 - INS 
 tpg|BK006946.2| 82391 + tpg|BK006946.2| 82052 - INS 
 tpg|BK006938.2| 480399 + tpg|BK006938.2| 480495 - INS 
 tpg|BK006938.2| 706224 + tpg|BK006938.2| 705828 - INS 
 tpg|BK006946.2| 483156 + tpg|BK006946.2| 483744 - INS 
 tpg|BK006946.2| 129053 + tpg|BK006946.2| 128602 - INS 
 tpg|BK006938.2| 932679 + tpg|BK006938.2| 932285 - INS 
 tpg|BK006946.2| 341493 + tpg|BK006946.2| 341876 - INS 
 tpg|BK006938.2| 1255482 + tpg|BK006938.2| 1255484 - INS 
 tpg|BK006938.2| 1026981 + tpg|BK006938.2| 1027402 - INS 
 tpg|BK006938.2| 19937 + tpg|BK006938.2| 19455 - INS 
 tpg|BK006938.2| 1021882 + tpg|BK006938.2| 1022155 - INS 
 tpg|BK006938.2| 120539 + tpg|BK006938.2| 120263 - INS 
 tpg|BK006938.2| 212404 + tpg|BK006938.2| 212186 - INS 
 tpg|BK006938.2| 335205 + tpg|BK006938.2| 334758 - INS 
 tpg|BK006946.2| 814279 + tpg|BK006946.2| 813565 - INS 
 tpg|BK006946.2| 705980 + tpg|BK006946.2| 705432 - INS 
 tpg|BK006938.2| 48832 + tpg|BK006938.2| 48192 - INS 
 tpg|BK006946.2| 915766 + tpg|BK006946.2| 916160 - INS 
 tpg|BK006946.2| 209985 + tpg|BK006946.2| 209692 - INS 
 tpg|BK006938.2| 1348859 + tpg|BK006938.2| 1348775 - INS 
 tpg|BK006946.2| 896424 + tpg|BK006946.2| 896606 - INS 
 tpg|BK006946.2| 33004 + tpg|BK006946.2| 32759 - INS 
 tpg|BK006946.2| 260179 + tpg|BK006946.2| 259671 - INS 
 tpg|BK006938.2| 456003 + tpg|BK006938.2| 455245 - INS 
 tpg|BK006946.2| 17239 + tpg|BK006946.2| 17405 - INS 
 tpg|BK006938.2| 381739 + tpg|BK006938.2| 381218 - INS 
 tpg|BK006938.2| 376400 + tpg|BK006938.2| 376327 - INS 
 tpg|BK006946.2| 536010 + tpg|BK006946.2| 535526 - INS 
 tpg|BK006938.2| 257231 + tpg|BK006938.2| 257451 - INS 
 tpg|BK006946.2| 529294 + tpg|BK006946.2| 529541 - INS 
 tpg|BK006946.2| 109732 + tpg|BK006946.2| 109626 - INS 
 tpg|BK006946.2| 842548 + tpg|BK006946.2| 842728 - INS 
 tpg|BK006946.2| 643763 + tpg|BK006946.2| 644099 - INS 
 tpg|BK006946.2| 629859 + tpg|BK006946.2| 629844 - INS 
 tpg|BK006946.2| 870153 + tpg|BK006946.2| 870011 - INS 
 tpg|BK006938.2| 1455899 + tpg|BK006938.2| 1456652 - INS 
 tpg|BK006946.2| 72304 + tpg|BK006946.2| 71996 - INS 
 tpg|BK006938.2| 527197 + tpg|BK006938.2| 527218 - INS 
 tpg|BK006938.2| 538521 + tpg|BK006938.2| 539227 - INS 
 tpg|BK006946.2| 400564 + tpg|BK006946.2| 399800 - INS 
 tpg|BK006938.2| 550358 + tpg|BK006938.2| 551026 - INS 
 tpg|BK006946.2| 848542 + tpg|BK006946.2| 848817 - INS 
 tpg|BK006938.2| 247688 + tpg|BK006938.2| 247308 - INS 
 tpg|BK006938.2| 520354 + tpg|BK006938.2| 520839 - INS 
 tpg|BK006946.2| 866312 + tpg|BK006946.2| 866327 - INS 
 tpg|BK006938.2| 1379558 + tpg|BK006938.2| 1380276 - INS 
 tpg|BK006938.2| 1356044 + tpg|BK006938.2| 1356348 - INS 
 tpg|BK006946.2| 291145 + tpg|BK006946.2| 291340 - INS 
 tpg|BK006938.2| 345037 + tpg|BK006938.2| 344598 - INS 
 tpg|BK006946.2| 237994 + tpg|BK006946.2| 237622 - INS 
 tpg|BK006938.2| 795126 + tpg|BK006938.2| 794604 - INS 
 tpg|BK006938.2| 1471646 + tpg|BK006938.2| 1471385 - INS 
 tpg|BK006938.2| 1337012 + tpg|BK006938.2| 1336505 - INS 
 tpg|BK006938.2| 748767 + tpg|BK006938.2| 748540 - INS 
 tpg|BK006946.2| 833479 + tpg|BK006946.2| 833992 - INS 
 tpg|BK006938.2| 791035 + tpg|BK006938.2| 790340 - INS 
 tpg|BK006938.2| 284622 + tpg|BK006938.2| 284979 - INS 
 tpg|BK006938.2| 780742 + tpg|BK006938.2| 780223 - INS 
 tpg|BK006946.2| 63664 + tpg|BK006946.2| 64030 - INS 
 tpg|BK006938.2| 782631 + tpg|BK006938.2| 782786 - INS 
 tpg|BK006938.2| 656327 + tpg|BK006938.2| 655625 - INS 
 tpg|BK006938.2| 785301 + tpg|BK006938.2| 785427 - INS 
 tpg|BK006938.2| 1517025 + tpg|BK006938.2| 1516722 - INS 
 tpg|BK006946.2| 592350 + tpg|BK006946.2| 591879 - INS 
 tpg|BK006938.2| 674511 + tpg|BK006938.2| 673899 - INS 
 tpg|BK006946.2| 779631 + tpg|BK006946.2| 779136 - INS 
 tpg|BK006938.2| 774772 + tpg|BK006938.2| 774532 - INS 
 tpg|BK006938.2| 227736 + tpg|BK006938.2| 228500 - INS 
 tpg|BK006938.2| 1503312 + tpg|BK006938.2| 1503238 - INS 
 tpg|BK006946.2| 367220 + tpg|BK006946.2| 367712 - INS 
 tpg|BK006938.2| 117531 + tpg|BK006938.2| 117445 - INS 
 tpg|BK006946.2| 20850 + tpg|BK006946.2| 20257 - INS 
 tpg|BK006938.2| 1499716 + tpg|BK006938.2| 1499582 - INS 
 tpg|BK006938.2| 1079945 + tpg|BK006938.2| 1079530 - INS 
 tpg|BK006938.2| 1484116 + tpg|BK006938.2| 1484105 - INS 
 tpg|BK006938.2| 1483483 + tpg|BK006938.2| 1482998 - INS 
 tpg|BK006946.2| 904079 + tpg|BK006946.2| 903958 - INS 
 tpg|BK006938.2| 1447781 + tpg|BK006938.2| 1447284 - INS 
 tpg|BK006946.2| 558192 + tpg|BK006946.2| 558160 - INS 
 tpg|BK006938.2| 710531 + tpg|BK006938.2| 710994 - INS 
 tpg|BK006938.2| 1422714 + tpg|BK006938.2| 1422244 - INS 
 tpg|BK006946.2| 203365 + tpg|BK006946.2| 203385 - INS 
 tpg|BK006938.2| 294782 + tpg|BK006938.2| 294851 - INS CTTTTTGCTC
 tpg|BK006938.2| 1121834 + tpg|BK006938.2| 1122031 - INS 
 tpg|BK006938.2| 187478 + tpg|BK006938.2| 187110 - INS 
 tpg|BK006938.2| 308344 + tpg|BK006938.2| 308869 - INS 
 tpg|BK006946.2| 573649 + tpg|BK006946.2| 573029 - INS 
 tpg|BK006938.2| 317584 + tpg|BK006938.2| 317026 - INS 
 tpg|BK006938.2| 902303 + tpg|BK006938.2| 902252 - INS 
 tpg|BK006938.2| 525619 + tpg|BK006938.2| 525221 - INS 
 tpg|BK006938.2| 156335 + tpg|BK006938.2| 155807 - INS 
 tpg|BK006938.2| 135054 + tpg|BK006938.2| 135457 - INS 
 tpg|BK006946.2| 888180 + tpg|BK006946.2| 887514 - INS 
 tpg|BK006938.2| 365022 + tpg|BK006938.2| 364436 - INS 
 tpg|BK006946.2| 307297 + tpg|BK006946.2| 306873 - INS 
 tpg|BK006938.2| 908816 + tpg|BK006938.2| 908508 - INS 
 tpg|BK006946.2| 154347 + tpg|BK006946.2| 154835 - INS 
 tpg|BK006938.2| 961646 + tpg|BK006938.2| 961903 - INS 
 tpg|BK006938.2| 970124 + tpg|BK006938.2| 970131 - INS 
 tpg|BK006938.2| 402243 + tpg|BK006938.2| 402875 - INS 
 tpg|BK006938.2| 405212 + tpg|BK006938.2| 405429 - INS GG
 tpg|BK006938.2| 58586 + tpg|BK006938.2| 58875 - INS 
 tpg|BK006938.2| 933295 + tpg|BK006938.2| 934033 - INS 
 tpg|BK006938.2| 608019 + tpg|BK006938.2| 608604 - INS 
 tpg|BK006938.2| 1234239 + tpg|BK006938.2| 1233635 - INS 
 tpg|BK006938.2| 1015561 + tpg|BK006938.2| 1015148 - INS 
 tpg|BK006938.2| 320312 + tpg|BK006938.2| 319970 - INS 
 tpg|BK006938.2| 1186107 + tpg|BK006938.2| 1186256 - INS 
 tpg|BK006938.2| 1176744 + tpg|BK006938.2| 1176315 - INS 
 tpg|BK006938.2| 378025 + tpg|BK006938.2| 377646 - INS 
 tpg|BK006938.2| 564263 + tpg|BK006938.2| 564375 - INS 
 tpg|BK006938.2| 488473 + tpg|BK006938.2| 488389 - INS 
 tpg|BK006938.2| 482975 + tpg|BK006938.2| 483271 - INS 
 tpg|BK006946.2| 862981 + tpg|BK006946.2| 862419 - INS 
 tpg|BK006938.2| 1163848 + tpg|BK006938.2| 1163506 - INS 
 tpg|BK006946.2| 424529 + tpg|BK006946.2| 424160 - INS 
 tpg|BK006938.2| 1332741 + tpg|BK006938.2| 1332319 - INS 
 tpg|BK006938.2| 526408 + tpg|BK006938.2| 525809 - INS 
 tpg|BK006946.2| 861397 + tpg|BK006946.2| 861197 - INS 
 tpg|BK006938.2| 1114158 + tpg|BK006938.2| 1113971 - INS 
 tpg|BK006938.2| 504656 + tpg|BK006938.2| 504072 - INS 
 tpg|BK006946.2| 627758 + tpg|BK006946.2| 627454 - INS 
 tpg|BK006938.2| 298867 + tpg|BK006938.2| 298942 - INS 
 tpg|BK006946.2| 85318 + tpg|BK006946.2| 85048 - INS 
 tpg|BK006938.2| 158376 + tpg|BK006938.2| 157981 - INS 
 tpg|BK006938.2| 275985 + tpg|BK006938.2| 275801 - INS 
 tpg|BK006938.2| 1181933 + tpg|BK006938.2| 1181321 - INS 
 tpg|BK006946.2| 109200 + tpg|BK006946.2| 108862 - INS 
 tpg|BK006938.2| 1228906 + tpg|BK006938.2| 1228313 - INS 
 tpg|BK006938.2| 1454608 + tpg|BK006938.2| 1453861 - INS 
 tpg|BK006946.2| 120589 + tpg|BK006946.2| 120576 - INS 
 tpg|BK006938.2| 310013 + tpg|BK006938.2| 309833 - INS 
 tpg|BK006938.2| 1167466 + tpg|BK006938.2| 1167076 - INS 
 tpg|BK006946.2| 645264 + tpg|BK006946.2| 644768 - INS 
 tpg|BK006946.2| 414128 + tpg|BK006946.2| 414879 - INS 
 tpg|BK006938.2| 476462 + tpg|BK006938.2| 476426 - INS 
 tpg|BK006946.2| 856453 + tpg|BK006946.2| 855717 - INS 
 tpg|BK006938.2| 100982 + tpg|BK006938.2| 101268 - INS 
 tpg|BK006938.2| 1220475 + tpg|BK006938.2| 1220013 - INS 
 tpg|BK006946.2| 635211 + tpg|BK006946.2| 635278 - INS 
 tpg|BK006938.2| 1381111 + tpg|BK006938.2| 1380762 - INS 
 tpg|BK006938.2| 684006 + tpg|BK006938.2| 684534 - INS 
 tpg|BK006938.2| 184955 + tpg|BK006938.2| 185219 - INS 
 tpg|BK006946.2| 425032 + tpg|BK006946.2| 425672 - INS 
 tpg|BK006938.2| 687683 + tpg|BK006938.2| 687486 - INS 
 tpg|BK006938.2| 1505505 + tpg|BK006938.2| 1505255 - INS 
 tpg|BK006946.2| 672991 + tpg|BK006946.2| 672639 - INS 
 tpg|BK006938.2| 79910 + tpg|BK006938.2| 79436 - INS 
 tpg|BK006938.2| 1235938 + tpg|BK006938.2| 1236486 - INS 
 tpg|BK006946.2| 417223 + tpg|BK006946.2| 416616 - INS 
 tpg|BK006938.2| 993918 + tpg|BK006938.2| 993542 - INS 
 tpg|BK006938.2| 1267945 + tpg|BK006938.2| 1268285 - INS 
 tpg|BK006938.2| 719714 + tpg|BK006938.2| 719843 - INS 
 tpg|BK006946.2| 69055 + tpg|BK006946.2| 69228 - INS 
 tpg|BK006946.2| 873424 + tpg|BK006946.2| 873235 - INS 
 tpg|BK006946.2| 889816 + tpg|BK006946.2| 889173 - INS 
 tpg|BK006938.2| 123270 + tpg|BK006938.2| 122503 - INS 
 tpg|BK006938.2| 1277329 + tpg|BK006938.2| 1276617 - INS 
 tpg|BK006946.2| 524294 + tpg|BK006946.2| 524988 - INS 
 tpg|BK006938.2| 1374299 + tpg|BK006938.2| 1373630 - INS 
 tpg|BK006946.2| 288289 + tpg|BK006946.2| 287838 - INS 
 tpg|BK006938.2| 818087 + tpg|BK006938.2| 817566 - INS GTAG
 tpg|BK006938.2| 1365616 + tpg|BK006938.2| 1365726 - INS 
 tpg|BK006946.2| 127485 + tpg|BK006946.2| 127339 - INS 
 tpg|BK006938.2| 763970 + tpg|BK006938.2| 764573 - INS 
 tpg|BK006938.2| 766333 + tpg|BK006938.2| 766736 - INS 
 tpg|BK006938.2| 339416 + tpg|BK006938.2| 339075 - INS 
 tpg|BK006946.2| 496948 + tpg|BK006946.2| 496525 - INS 
 tpg|BK006946.2| 510355 + tpg|BK006946.2| 509845 - INS 
 tpg|BK006946.2| 119638 + tpg|BK006946.2| 119703 - INS 
 tpg|BK006938.2| 916961 + tpg|BK006938.2| 916639 - INS 
 tpg|BK006938.2| 76016 + tpg|BK006938.2| 75402 - INS 
 tpg|BK006938.2| 943818 + tpg|BK006938.2| 943615 - INS 
 tpg|BK006938.2| 448292 + tpg|BK006938.2| 448329 - INS 
 tpg|BK006938.2| 404513 + tpg|BK006938.2| 404267 - INS 
 tpg|BK006938.2| 471915 + tpg|BK006938.2| 471372 - INS 
 tpg|BK006946.2| 285741 + tpg|BK006946.2| 286106 - INS 
 tpg|BK006938.2| 1304303 + tpg|BK006938.2| 1304971 - INS 
 tpg|BK006938.2| 739945 + tpg|BK006938.2| 739440 - INS 
 tpg|BK006938.2| 605804 + tpg|BK006938.2| 605892 - INS 
 tpg|BK006938.2| 819441 + tpg|BK006938.2| 818825 - INS 
 tpg|BK006938.2| 1149946 + tpg|BK006938.2| 1149743 - INS 
 tpg|BK006938.2| 689835 + tpg|BK006938.2| 690342 - INS 
 tpg|BK006946.2| 449850 + tpg|BK006946.2| 449999 - INS 
 tpg|BK006938.2| 32148 + tpg|BK006938.2| 32771 - INS 
 tpg|BK006946.2| 469923 + tpg|BK006946.2| 470032 - INS 
 tpg|BK006938.2| 51341 + tpg|BK006938.2| 51315 - INS 
 tpg|BK006938.2| 667798 + tpg|BK006938.2| 667685 - INS 
 tpg|BK006946.2| 549663 + tpg|BK006946.2| 550250 - INS 
 tpg|BK006946.2| 546973 + tpg|BK006946.2| 546929 - INS 
 tpg|BK006946.2| 519031 + tpg|BK006946.2| 519306 - INS 
 tpg|BK006938.2| 1026186 + tpg|BK006938.2| 1025663 - INS 
 tpg|BK006938.2| 341574 + tpg|BK006938.2| 341824 - INS 
 tpg|BK006946.2| 769601 + tpg|BK006946.2| 770287 - INS 
 tpg|BK006946.2| 534808 + tpg|BK006946.2| 534798 - INS 
 tpg|BK006946.2| 546007 + tpg|BK006946.2| 545617 - INS 
 tpg|BK006938.2| 812100 + tpg|BK006938.2| 811680 - INS 
 tpg|BK006946.2| 291604 + tpg|BK006946.2| 292249 - INS 
 tpg|BK006938.2| 751714 + tpg|BK006938.2| 751317 - INS 
 tpg|BK006938.2| 823513 + tpg|BK006938.2| 823324 - INS 
 tpg|BK006946.2| 578109 + tpg|BK006946.2| 577752 - INS 
 tpg|BK006938.2| 222397 + tpg|BK006938.2| 221623 - INS 
 tpg|BK006946.2| 787629 + tpg|BK006946.2| 786862 - INS 
 tpg|BK006938.2| 1511466 + tpg|BK006938.2| 1511207 - INS 
 tpg|BK006938.2| 803607 + tpg|BK006938.2| 803205 - INS 
 tpg|BK006938.2| 765430 + tpg|BK006938.2| 765245 - INS 
 tpg|BK006946.2| 722270 + tpg|BK006946.2| 722504 - INS 
 tpg|BK006938.2| 1151437 + tpg|BK006938.2| 1150917 - INS 
 tpg|BK006946.2| 168414 + tpg|BK006946.2| 167889 - INS 
 tpg|BK006938.2| 50158 + tpg|BK006938.2| 49771 - INS 
 tpg|BK006938.2| 1316645 + tpg|BK006938.2| 1316608 - INS 
 tpg|BK006946.2| 62728 + tpg|BK006946.2| 62740 - INS 
 tpg|BK006938.2| 1342807 + tpg|BK006938.2| 1342895 - INS 
 tpg|BK006938.2| 405873 + tpg|BK006938.2| 406300 - INS 
 tpg|BK006938.2| 1112219 + tpg|BK006938.2| 1112173 - INS 
 tpg|BK006946.2| 381378 + tpg|BK006946.2| 381278 - INS 
 tpg|BK006938.2| 1289563 + tpg|BK006938.2| 1289628 - INS 
 tpg|BK006946.2| 812442 + tpg|BK006946.2| 812824 - INS 
 tpg|BK006938.2| 362407 + tpg|BK006938.2| 362145 - INS 
 tpg|BK006938.2| 949928 + tpg|BK006938.2| 949602 - INS 
 tpg|BK006938.2| 592090 + tpg|BK006938.2| 591610 - INS 
 tpg|BK006946.2| 329196 + tpg|BK006946.2| 328537 - INS 
 tpg|BK006938.2| 602810 + tpg|BK006938.2| 602248 - INS 
 tpg|BK006938.2| 224510 + tpg|BK006938.2| 224233 - INS 
 tpg|BK006946.2| 703860 + tpg|BK006946.2| 703522 - INS 
 tpg|BK006938.2| 496533 + tpg|BK006938.2| 495994 - INS 
 tpg|BK006938.2| 901461 + tpg|BK006938.2| 901512 - INS 
 tpg|BK006946.2| 320881 + tpg|BK006946.2| 320165 - INS 
 tpg|BK006938.2| 825821 + tpg|BK006938.2| 826365 - INS 
 tpg|BK006938.2| 1102980 + tpg|BK006938.2| 1102565 - INS 
 tpg|BK006946.2| 652190 + tpg|BK006946.2| 651917 - INS 
 tpg|BK006938.2| 1243062 + tpg|BK006938.2| 1242641 - INS 
 tpg|BK006946.2| 650429 + tpg|BK006946.2| 650671 - INS 
 tpg|BK006938.2| 1024801 + tpg|BK006938.2| 1024437 - INS 
 tpg|BK006938.2| 1200324 + tpg|BK006938.2| 1199794 - INS 
 tpg|BK006938.2| 374846 + tpg|BK006938.2| 374655 - INS 
 tpg|BK006946.2| 144681 + tpg|BK006946.2| 145082 - INS 
 tpg|BK006938.2| 425323 + tpg|BK006938.2| 424646 - INS 
 tpg|BK006938.2| 709910 + tpg|BK006938.2| 710013 - INS 
 tpg|BK006946.2| 801262 + tpg|BK006946.2| 801630 - INS 
 tpg|BK006938.2| 1224882 + tpg|BK006938.2| 1224837 - INS 
 tpg|BK006938.2| 387309 + tpg|BK006938.2| 387502 - INS 
 tpg|BK006946.2| 824239 + tpg|BK006946.2| 823544 - INS 
 tpg|BK006946.2| 636532 + tpg|BK006946.2| 636678 - INS 
 tpg|BK006946.2| 355906 + tpg|BK006946.2| 356610 - INS 
 tpg|BK006938.2| 255761 + tpg|BK006938.2| 256002 - INS 
 tpg|BK006938.2| 580332 + tpg|BK006938.2| 580011 - INS 
 tpg|BK006946.2| 859053 + tpg|BK006946.2| 859648 - INS 
 tpg|BK006938.2| 1229595 + tpg|BK006938.2| 1229156 - INS 
 tpg|BK006938.2| 972501 + tpg|BK006938.2| 972241 - INS 
 tpg|BK006938.2| 666712 + tpg|BK006938.2| 666218 - INS 
 tpg|BK006946.2| 300374 + tpg|BK006946.2| 299959 - INS 
 tpg|BK006938.2| 1206168 + tpg|BK006938.2| 1206505 - INS 
 tpg|BK006938.2| 1010339 + tpg|BK006938.2| 1010743 - INS 
 tpg|BK006946.2| 522621 + tpg|BK006946.2| 523290 - INS 
 tpg|BK006938.2| 58166 + tpg|BK006938.2| 57632 - INS 
 tpg|BK006946.2| 77967 + tpg|BK006946.2| 78403 - INS 
 tpg|BK006946.2| 428216 + tpg|BK006946.2| 428119 - INS 
 tpg|BK006938.2| 74487 + tpg|BK006938.2| 74069 - INS 
 tpg|BK006938.2| 1162389 + tpg|BK006938.2| 1161819 - INS 
 tpg|BK006938.2| 814187 + tpg|BK006938.2| 813993 - INS 
 tpg|BK006946.2| 428899 + tpg|BK006946.2| 428759 - INS 
 tpg|BK006938.2| 1349349 + tpg|BK006938.2| 1349844 - INS 
 tpg|BK006938.2| 824722 + tpg|BK006938.2| 824460 - INS 
 tpg|BK006938.2| 1409277 + tpg|BK006938.2| 1409369 - INS 
 tpg|BK006946.2| 726899 + tpg|BK006946.2| 727231 - INS 
 tpg|BK006938.2| 324313 + tpg|BK006938.2| 323969 - INS 
 tpg|BK006938.2| 917445 + tpg|BK006938.2| 917700 - INS 
 tpg|BK006938.2| 979644 + tpg|BK006938.2| 979169 - INS 
 tpg|BK006946.2| 785459 + tpg|BK006946.2| 785810 - INS 
 tpg|BK006938.2| 1421290 + tpg|BK006938.2| 1421589 - INS 
 tpg|BK006938.2| 1028524 + tpg|BK006938.2| 1029054 - INS 
 tpg|BK006938.2| 69407 + tpg|BK006938.2| 68983 - INS 
 tpg|BK006946.2| 143524 + tpg|BK006946.2| 142780 - INS 
 tpg|BK006938.2| 323707 + tpg|BK006938.2| 323170 - INS 
 tpg|BK006938.2| 1267114 + tpg|BK006938.2| 1266943 - INS 
 tpg|BK006946.2| 97509 + tpg|BK006946.2| 97896 - INS 
 tpg|BK006938.2| 1015034 + tpg|BK006938.2| 1014699 - INS 
 tpg|BK006938.2| 191528 + tpg|BK006938.2| 191476 - INS 
 tpg|BK006946.2| 296990 + tpg|BK006946.2| 296323 - INS 
 tpg|BK006938.2| 959370 + tpg|BK006938.2| 959185 - INS 
 tpg|BK006946.2| 803928 + tpg|BK006946.2| 803256 - INS 
 tpg|BK006938.2| 846602 + tpg|BK006938.2| 846473 - INS 
 tpg|BK006946.2| 708764 + tpg|BK006946.2| 708347 - INS 
 tpg|BK006946.2| 65956 + tpg|BK006946.2| 66508 - INS 
 tpg|BK006938.2| 699778 + tpg|BK006938.2| 699587 - INS 
 tpg|BK006938.2| 1128756 + tpg|BK006938.2| 1128175 - INS 
 tpg|BK006938.2| 280820 + tpg|BK006938.2| 280341 - INS 
 tpg|BK006938.2| 865186 + tpg|BK006938.2| 865635 - INS 
 tpg|BK006938.2| 849620 + tpg|BK006938.2| 849324 - INS 
 tpg|BK006938.2| 286914 + tpg|BK006938.2| 286219 - INS 
 tpg|BK006938.2| 558796 + tpg|BK006938.2| 559434 - INS 
 tpg|BK006938.2| 1202123 + tpg|BK006938.2| 1201768 - INS 
 tpg|BK006938.2| 1103542 + tpg|BK006938.2| 1104014 - INS 
 tpg|BK006938.2| 1133749 + tpg|BK006938.2| 1133319 - INS 
 tpg|BK006938.2| 254980 + tpg|BK006938.2| 254965 - INS 
 tpg|BK006938.2| 81976 + tpg|BK006938.2| 81430 - INS 
 tpg|BK006938.2| 1245960 + tpg|BK006938.2| 1246597 - INS 
 tpg|BK006938.2| 1457075 + tpg|BK006938.2| 1457801 - INS 
 tpg|BK006938.2| 892528 + tpg|BK006938.2| 891798 - INS 
 tpg|BK006938.2| 1465112 + tpg|BK006938.2| 1464933 - INS 
 tpg|BK006946.2| 891831 + tpg|BK006946.2| 892118 - INS 
 tpg|BK006938.2| 586998 + tpg|BK006938.2| 586812 - INS 
 tpg|BK006938.2| 427412 + tpg|BK006938.2| 426716 - INS 
 tpg|BK006938.2| 1039474 + tpg|BK006938.2| 1039207 - INS 
 tpg|BK006938.2| 1342322 + tpg|BK006938.2| 1341594 - INS 
 tpg|BK006938.2| 670916 + tpg|BK006938.2| 670641 - INS 
 tpg|BK006938.2| 277271 + tpg|BK006938.2| 276853 - INS 
 tpg|BK006938.2| 249020 + tpg|BK006938.2| 248381 - INS 
 tpg|BK006938.2| 1303103 + tpg|BK006938.2| 1302800 - INS 
 tpg|BK006938.2| 1334476 + tpg|BK006938.2| 1333809 - INS 
 tpg|BK006938.2| 466991 + tpg|BK006938.2| 466663 - INS 
 tpg|BK006938.2| 1224157 + tpg|BK006938.2| 1224013 - INS 
 tpg|BK006938.2| 139979 + tpg|BK006938.2| 140177 - INS 
 tpg|BK006938.2| 111849 + tpg|BK006938.2| 111775 - INS 
 tpg|BK006938.2| 513369 + tpg|BK006938.2| 512805 - INS 
 tpg|BK006938.2| 1235231 + tpg|BK006938.2| 1234772 - INS 
 tpg|BK006938.2| 432995 + tpg|BK006938.2| 432306 - INS 
 tpg|BK006938.2| 720862 + tpg|BK006938.2| 721128 - INS 
 tpg|BK006938.2| 1217911 + tpg|BK006938.2| 1217819 - INS 
 tpg|BK006938.2| 1201001 + tpg|BK006938.2| 1201188 - INS 
 tpg|BK006938.2| 1321453 + tpg|BK006938.2| 1321198 - INS 
 tpg|BK006938.2| 1263117 + tpg|BK006938.2| 1263214 - INS 
 tpg|BK006938.2| 857323 + tpg|BK006938.2| 857230 - INS 
 tpg|BK006938.2| 995256 + tpg|BK006938.2| 995165 - INS 
 tpg|BK006938.2| 899510 + tpg|BK006938.2| 898881 - INS 
 tpg|BK006938.2| 583314 + tpg|BK006938.2| 583626 - INS 
 tpg|BK006938.2| 896220 + tpg|BK006938.2| 895812 - INS 
 tpg|BK006938.2| 1371505 + tpg|BK006938.2| 1371202 - INS 
 tpg|BK006938.2| 167332 + tpg|BK006938.2| 167582 - INS 
 tpg|BK006946.2| 382714 + tpg|BK006946.2| 382348 - INS 
 tpg|BK006938.2| 24673 + tpg|BK006938.2| 24735 - INS 
 tpg|BK006938.2| 161418 + tpg|BK006938.2| 160889 - INS 
 tpg|BK006938.2| 424281 + tpg|BK006938.2| 424160 - INS 
 tpg|BK006938.2| 1325717 + tpg|BK006938.2| 1325477 - INS 
 tpg|BK006946.2| 288841 + tpg|BK006946.2| 288962 - INS 
 tpg|BK006938.2| 1482142 + tpg|BK006938.2| 1482456 - INS 
 tpg|BK006938.2| 386482 + tpg|BK006938.2| 385834 - INS 
 tpg|BK006938.2| 1487644 + tpg|BK006938.2| 1487079 - INS 
 tpg|BK006938.2| 966533 + tpg|BK006938.2| 966097 - INS 
 tpg|BK006946.2| 565938 + tpg|BK006946.2| 565813 - INS 
 tpg|BK006938.2| 834488 + tpg|BK006938.2| 834544 - INS 
 tpg|BK006938.2| 872194 + tpg|BK006938.2| 871773 - INS 
 tpg|BK006938.2| 808381 + tpg|BK006938.2| 808172 - INS 
 tpg|BK006938.2| 1134299 + tpg|BK006938.2| 1133736 - INS 
 tpg|BK006946.2| 205207 + tpg|BK006946.2| 204518 - INS 
 tpg|BK006938.2| 17549 + tpg|BK006938.2| 18098 - INS 
 tpg|BK006938.2| 1159729 + tpg|BK006938.2| 1159410 - INS 
 tpg|BK006938.2| 1501881 + tpg|BK006938.2| 1501403 - INS 
 tpg|BK006938.2| 345438 + tpg|BK006938.2| 345405 - INS 
 tpg|BK006946.2| 667182 + tpg|BK006946.2| 666557 - INS 
 tpg|BK006938.2| 119189 + tpg|BK006938.2| 119700 - INS 
 tpg|BK006938.2| 747114 + tpg|BK006938.2| 746816 - INS 
 tpg|BK006946.2| 839625 + tpg|BK006946.2| 840089 - INS 
 tpg|BK006946.2| 129683 + tpg|BK006946.2| 129242 - INS 
 tpg|BK006938.2| 1418116 + tpg|BK006938.2| 1418191 - INS 
 tpg|BK006946.2| 876211 + tpg|BK006946.2| 875946 - INS 
 tpg|BK006938.2| 370324 + tpg|BK006938.2| 370020 - INS 
 tpg|BK006938.2| 412710 + tpg|BK006938.2| 413187 - INS 
 tpg|BK006946.2| 413621 + tpg|BK006946.2| 413317 - INS 
 tpg|BK006938.2| 437533 + tpg|BK006938.2| 437978 - INS 
 tpg|BK006938.2| 327690 + tpg|BK006938.2| 327471 - INS 
 tpg|BK006946.2| 294803 + tpg|BK006946.2| 294531 - INS 
 tpg|BK006938.2| 713046 + tpg|BK006938.2| 712448 - INS 
 tpg|BK006938.2| 512857 + tpg|BK006938.2| 512405 - INS 
 tpg|BK006938.2| 576635 + tpg|BK006938.2| 576474 - INS 
 tpg|BK006946.2| 195747 + tpg|BK006946.2| 196213 - INS 
 tpg|BK006938.2| 313064 + tpg|BK006938.2| 312496 - INS 
 tpg|BK006938.2| 326222 + tpg|BK006938.2| 326232 - INS 
 tpg|BK006938.2| 118574 + tpg|BK006938.2| 118390 - INS 
 tpg|BK006938.2| 1326499 + tpg|BK006938.2| 1326220 - INS 
 tpg|BK006938.2| 555637 + tpg|BK006938.2| 555628 - INS 
 tpg|BK006938.2| 428312 + tpg|BK006938.2| 427720 - INS 
 tpg|BK006938.2| 442553 + tpg|BK006938.2| 442241 - INS 
 tpg|BK006938.2| 987638 + tpg|BK006938.2| 987058 - INS 
 tpg|BK006938.2| 626905 + tpg|BK006938.2| 626215 - INS 
 tpg|BK006946.2| 354649 + tpg|BK006946.2| 355077 - INS 
 tpg|BK006938.2| 365401 + tpg|BK006938.2| 365093 - INS 
 tpg|BK006938.2| 180118 + tpg|BK006938.2| 179612 - INS 
 tpg|BK006938.2| 457843 + tpg|BK006938.2| 458286 - INS 
 tpg|BK006946.2| 913512 + tpg|BK006946.2| 913629 - INS 
 tpg|BK006938.2| 1028202 + tpg|BK006938.2| 1028690 - INS 
 tpg|BK006946.2| 844598 + tpg|BK006946.2| 843953 - INS 
 tpg|BK006938.2| 1121172 + tpg|BK006938.2| 1120971 - INS 
 tpg|BK006938.2| 144099 + tpg|BK006938.2| 143775 - INS 
 tpg|BK006946.2| 242564 + tpg|BK006946.2| 242512 - INS 
 tpg|BK006938.2| 811444 + tpg|BK006938.2| 811231 - INS 
 tpg|BK006938.2| 504056 + tpg|BK006938.2| 503591 - INS 
 tpg|BK006946.2| 851741 + tpg|BK006946.2| 851860 - INS 
 tpg|BK006938.2| 1333185 + tpg|BK006938.2| 1332971 - INS 
 tpg|BK006938.2| 892918 + tpg|BK006938.2| 892788 - INS 
 tpg|BK006946.2| 483765 + tpg|BK006946.2| 484305 - INS 
 tpg|BK006938.2| 822541 + tpg|BK006938.2| 821963 - INS 
 tpg|BK006938.2| 439200 + tpg|BK006938.2| 439089 - INS 
 tpg|BK006938.2| 335581 + tpg|BK006938.2| 335716 - INS 
 tpg|BK006938.2| 510090 + tpg|BK006938.2| 509338 - INS 
 tpg|BK006938.2| 401527 + tpg|BK006938.2| 401382 - INS 
 tpg|BK006938.2| 960422 + tpg|BK006938.2| 959802 - INS 
 tpg|BK006946.2| 537250 + tpg|BK006946.2| 536865 - INS 
 tpg|BK006938.2| 286187 + tpg|BK006938.2| 285690 - INS 
 tpg|BK006946.2| 526578 + tpg|BK006946.2| 526193 - INS 
 tpg|BK006938.2| 624583 + tpg|BK006938.2| 624229 - INS 
 tpg|BK006938.2| 323062 + tpg|BK006938.2| 322496 - INS 
 tpg|BK006946.2| 781688 + tpg|BK006946.2| 781415 - INS 
 tpg|BK006938.2| 475039 + tpg|BK006938.2| 474778 - INS 
 tpg|BK006938.2| 1512910 + tpg|BK006938.2| 1513608 - INS 
 tpg|BK006938.2| 563421 + tpg|BK006938.2| 562948 - INS 
 tpg|BK006938.2| 1462453 + tpg|BK006938.2| 1461892 - INS 
 tpg|BK006946.2| 433041 + tpg|BK006946.2| 432778 - INS 
 tpg|BK006938.2| 1346829 + tpg|BK006938.2| 1347150 - INS 
 tpg|BK006938.2| 1352649 + tpg|BK006938.2| 1352165 - INS 
 tpg|BK006938.2| 679278 + tpg|BK006938.2| 679169 - INS 
 tpg|BK006946.2| 193412 + tpg|BK006946.2| 193230 - INS 
 tpg|BK006938.2| 519702 + tpg|BK006938.2| 519293 - INS 
 tpg|BK006938.2| 1488271 + tpg|BK006938.2| 1487736 - INS 
 tpg|BK006938.2| 973017 + tpg|BK006938.2| 973083 - INS 
 tpg|BK006938.2| 354477 + tpg|BK006938.2| 354468 - INS 
 tpg|BK006946.2| 473251 + tpg|BK006946.2| 472992 - INS 
 tpg|BK006938.2| 951914 + tpg|BK006938.2| 951874 - INS 
 tpg|BK006938.2| 1197157 + tpg|BK006938.2| 1196702 - INS 
 tpg|BK006938.2| 70056 + tpg|BK006938.2| 69667 - INS 
 tpg|BK006946.2| 251207 + tpg|BK006946.2| 251365 - INS 
 tpg|BK006938.2| 208006 + tpg|BK006938.2| 207795 - INS 
 tpg|BK006938.2| 1202666 + tpg|BK006938.2| 1203292 - INS 
 tpg|BK006946.2| 590826 + tpg|BK006946.2| 590794 - INS 
 tpg|BK006938.2| 433700 + tpg|BK006938.2| 433599 - INS 
 tpg|BK006946.2| 460314 + tpg|BK006946.2| 460990 - INS 
 tpg|BK006938.2| 752519 + tpg|BK006938.2| 752054 - INS 
 tpg|BK006938.2| 1320828 + tpg|BK006938.2| 1320347 - INS 
 tpg|BK006938.2| 961073 + tpg|BK006938.2| 961212 - INS 
 tpg|BK006946.2| 453193 + tpg|BK006946.2| 452575 - INS 
 tpg|BK006938.2| 45506 + tpg|BK006938.2| 45295 - INS 
 tpg|BK006938.2| 1424798 + tpg|BK006938.2| 1424516 - INS 
 tpg|BK006946.2| 589165 + tpg|BK006946.2| 588476 - INS 
 tpg|BK006946.2| 879993 + tpg|BK006946.2| 879673 - INS 
 tpg|BK006946.2| 309922 + tpg|BK006946.2| 309677 - INS 
 tpg|BK006946.2| 879061 + tpg|BK006946.2| 878840 - INS 
 tpg|BK006946.2| 439379 + tpg|BK006946.2| 439015 - INS 
 tpg|BK006946.2| 58719 + tpg|BK006946.2| 58897 - INS 
 tpg|BK006946.2| 618961 + tpg|BK006946.2| 619103 - INS 
 tpg|BK006946.2| 788457 + tpg|BK006946.2| 788408 - INS 
 tpg|BK006946.2| 157748 + tpg|BK006946.2| 158389 - INS 
 tpg|BK006946.2| 799246 + tpg|BK006946.2| 798594 - INS 
 tpg|BK006946.2| 631413 + tpg|BK006946.2| 632085 - INS 
 tpg|BK006946.2| 152463 + tpg|BK006946.2| 152333 - INS 
 tpg|BK006946.2| 303022 + tpg|BK006946.2| 303343 - INS 
 tpg|BK006946.2| 342533 + tpg|BK006946.2| 342701 - INS 
 tpg|BK006946.2| 105707 + tpg|BK006946.2| 105410 - INS 
 tpg|BK006946.2| 701361 + tpg|BK006946.2| 701525 - INS 
 tpg|BK006946.2| 675716 + tpg|BK006946.2| 675266 - INS 
 tpg|BK006946.2| 638043 + tpg|BK006946.2| 637491 - INS 
 tpg|BK006946.2| 93905 + tpg|BK006946.2| 94125 - INS 
 tpg|BK006946.2| 395584 + tpg|BK006946.2| 395244 - INS 
 tpg|BK006946.2| 847016 + tpg|BK006946.2| 847188 - INS 
 tpg|BK006946.2| 840503 + tpg|BK006946.2| 840965 - INS 
 tpg|BK006946.2| 620378 + tpg|BK006946.2| 620616 - INS 
 tpg|BK006946.2| 436440 + tpg|BK006946.2| 436272 - INS 
 tpg|BK006946.2| 57679 + tpg|BK006946.2| 57475 - INS 
 tpg|BK006946.2| 458655 + tpg|BK006946.2| 457985 - INS 
 tpg|BK006946.2| 695458 + tpg|BK006946.2| 695480 - INS 
 tpg|BK006946.2| 36169 + tpg|BK006946.2| 36021 - INS 
 tpg|BK006946.2| 22968 + tpg|BK006946.2| 22690 - INS 
 tpg|BK006946.2| 598488 + tpg|BK006946.2| 598066 - INS 
 tpg|BK006946.2| 457081 + tpg|BK006946.2| 457187 - INS 
 tpg|BK006946.2| 906233 + tpg|BK006946.2| 905966 - INS 
 tpg|BK006946.2| 245496 + tpg|BK006946.2| 244818 - INS GTA
 tpg|BK006946.2| 756662 + tpg|BK006946.2| 756445 - INS 
 tpg|BK006946.2| 685647 + tpg|BK006946.2| 685204 - INS 
 tpg|BK006946.2| 816718 + tpg|BK006946.2| 816669 - INS 
 tpg|BK006946.2| 521939 + tpg|BK006946.2| 522134 - INS 
 tpg|BK006946.2| 162699 + tpg|BK006946.2| 162667 - INS 
 tpg|BK006946.2| 645764 + tpg|BK006946.2| 645628 - INS 
 tpg|BK006946.2| 298236 + tpg|BK006946.2| 298024 - INS 
 tpg|BK006946.2| 73837 + tpg|BK006946.2| 74057 - INS 
 tpg|BK006946.2| 615338 + tpg|BK006946.2| 615312 - INS 
 tpg|BK006946.2| 165603 + tpg|BK006946.2| 165245 - INS 
 tpg|BK006946.2| 77500 + tpg|BK006946.2| 77846 - INS 
 tpg|BK006946.2| 92383 + tpg|BK006946.2| 92583 - INS 
 tpg|BK006946.2| 476706 + tpg|BK006946.2| 476995 - INS 
 tpg|BK006946.2| 541038 + tpg|BK006946.2| 541343 - INS 
 tpg|BK006946.2| 23791 + tpg|BK006946.2| 23605 - INS 
 tpg|BK006946.2| 542338 + tpg|BK006946.2| 541793 - INS 
 tpg|BK006946.2| 446411 + tpg|BK006946.2| 446664 - INS 
 tpg|BK006946.2| 491021 + tpg|BK006946.2| 491215 - INS 
 tpg|BK006946.2| 912094 + tpg|BK006946.2| 911862 - INS 
 tpg|BK006946.2| 821206 + tpg|BK006946.2| 821906 - INS GGGAA
 tpg|BK006946.2| 471389 + tpg|BK006946.2| 472015 - INS 
 tpg|BK006946.2| 579112 + tpg|BK006946.2| 579767 - INS 
 tpg|BK006946.2| 444006 + tpg|BK006946.2| 443264 - INS 
 tpg|BK006946.2| 726322 + tpg|BK006946.2| 725758 - INS 
 tpg|BK006946.2| 758183 + tpg|BK006946.2| 757922 - INS 
 tpg|BK006946.2| 676502 + tpg|BK006946.2| 676194 - INS 
 tpg|BK006946.2| 854338 + tpg|BK006946.2| 855094 - INS 
 tpg|BK006946.2| 141801 + tpg|BK006946.2| 141368 - INS 
 tpg|BK006946.2| 427322 + tpg|BK006946.2| 426911 - INS 
 tpg|BK006946.2| 430788 + tpg|BK006946.2| 430512 - INS 
 tpg|BK006946.2| 163410 + tpg|BK006946.2| 163774 - INS 
 tpg|BK006946.2| 171334 + tpg|BK006946.2| 171431 - INS 
 tpg|BK006946.2| 791574 + tpg|BK006946.2| 791422 - INS 
 tpg|BK006946.2| 469156 + tpg|BK006946.2| 468711 - INS 
 tpg|BK006946.2| 574465 + tpg|BK006946.2| 574049 - INS 
 tpg|BK006946.2| 40589 + tpg|BK006946.2| 40882 - INS 
 tpg|BK006946.2| 482205 + tpg|BK006946.2| 482125 - INS 
 tpg|BK006946.2| 740469 + tpg|BK006946.2| 741222 - INS 
 tpg|BK006946.2| 742196 + tpg|BK006946.2| 742339 - INS 
 tpg|BK006946.2| 233268 + tpg|BK006946.2| 232898 - INS 
 tpg|BK006946.2| 227599 + tpg|BK006946.2| 226849 - INS 
 tpg|BK006946.2| 248830 + tpg|BK006946.2| 249157 - INS 
 tpg|BK006946.2| 508381 + tpg|BK006946.2| 508585 - INS 
 tpg|BK006946.2| 912885 + tpg|BK006946.2| 912599 - INS 
 tpg|BK006946.2| 217632 + tpg|BK006946.2| 218187 - INS 
 tpg|BK006946.2| 213035 + tpg|BK006946.2| 212566 - INS 
 tpg|BK006946.2| 783378 + tpg|BK006946.2| 782605 - INS 
 tpg|BK006946.2| 24642 + tpg|BK006946.2| 24878 - INS 
 tpg|BK006946.2| 283405 + tpg|BK006946.2| 282799 - INS GCTGC
 tpg|BK006946.2| 604178 + tpg|BK006946.2| 603998 - INS 
 tpg|BK006946.2| 161585 + tpg|BK006946.2| 161217 - INS 
 tpg|BK006946.2| 804560 + tpg|BK006946.2| 803971 - INS 
 tpg|BK006946.2| 76619 + tpg|BK006946.2| 76712 - INS 
 tpg|BK006946.2| 697945 + tpg|BK006946.2| 697562 - INS 
 tpg|BK006946.2| 420134 + tpg|BK006946.2| 420282 - INS 
 tpg|BK006946.2| 858202 + tpg|BK006946.2| 857911 - INS 
 tpg|BK006946.2| 853674 + tpg|BK006946.2| 853349 - INS 
 tpg|BK006946.2| 95937 + tpg|BK006946.2| 96100 - INS 
 tpg|BK006946.2| 669102 + tpg|BK006946.2| 669404 - INS 
 tpg|BK006946.2| 668274 + tpg|BK006946.2| 667744 - INS 
 tpg|BK006946.2| 830782 + tpg|BK006946.2| 830632 - INS 
 tpg|BK006946.2| 391470 + tpg|BK006946.2| 390888 - INS 
 tpg|BK006946.2| 380288 + tpg|BK006946.2| 380354 - INS 
 tpg|BK006946.2| 113489 + tpg|BK006946.2| 112850 - INS 
 tpg|BK006946.2| 653060 + tpg|BK006946.2| 652621 - INS 
 tpg|BK006946.2| 396861 + tpg|BK006946.2| 396505 - INS 
 tpg|BK006946.2| 50710 + tpg|BK006946.2| 50461 - INS 
 tpg|BK006946.2| 904837 + tpg|BK006946.2| 904542 - INS 
 tpg|BK006946.2| 730385 + tpg|BK006946.2| 730084 - INS 
 tpg|BK006946.2| 761910 + tpg|BK006946.2| 761649 - INS 
 tpg|BK006946.2| 681163 + tpg|BK006946.2| 681879 - INS 
 tpg|BK006946.2| 829725 + tpg|BK006946.2| 829324 - INS 
 tpg|BK006946.2| 605268 + tpg|BK006946.2| 605995 - INS 
 tpg|BK006946.2| 117327 + tpg|BK006946.2| 116620 - INS 
 tpg|BK006946.2| 282030 + tpg|BK006946.2| 282012 - INS 
 tpg|BK006946.2| 123664 + tpg|BK006946.2| 123483 - INS 
 tpg|BK006946.2| 626640 + tpg|BK006946.2| 626014 - INS 
 tpg|BK006946.2| 809654 + tpg|BK006946.2| 809211 - INS 
 tpg|BK006946.2| 314760 + tpg|BK006946.2| 315299 - INS 
 tpg|BK006946.2| 384824 + tpg|BK006946.2| 384063 - INS 
 tpg|BK006946.2| 99408 + tpg|BK006946.2| 99049 - INS 
 tpg|BK006946.2| 789283 + tpg|BK006946.2| 788825 - INS 
 tpg|BK006946.2| 506439 + tpg|BK006946.2| 506983 - INS 
 tpg|BK006946.2| 191577 + tpg|BK006946.2| 192054 - INS 
 tpg|BK006946.2| 139002 + tpg|BK006946.2| 138480 - INS 
 tpg|BK006946.2| 678132 + tpg|BK006946.2| 677484 - INS 
 tpg|BK006946.2| 330671 + tpg|BK006946.2| 330113 - INS 
 tpg|BK006946.2| 70989 + tpg|BK006946.2| 70530 - INS 
 tpg|BK006946.2| 490094 + tpg|BK006946.2| 490247 - INS 
 tpg|BK006946.2| 277064 + tpg|BK006946.2| 276835 - INS 
 tpg|BK006946.2| 21740 + tpg|BK006946.2| 21791 - INS 
 tpg|BK006946.2| 246749 + tpg|BK006946.2| 246857 - INS 
 tpg|BK006946.2| 379280 + tpg|BK006946.2| 378513 - INS 
 tpg|BK006946.2| 401635 + tpg|BK006946.2| 401028 - INS 
 tpg|BK006946.2| 385920 + tpg|BK006946.2| 386326 - INS 
 tpg|BK006946.2| 131383 + tpg|BK006946.2| 131264 - INS 
 tpg|BK006946.2| 792611 + tpg|BK006946.2| 792810 - INS 
 tpg|BK006946.2| 569376 + tpg|BK006946.2| 570143 - INS 
 tpg|BK006946.2| 322735 + tpg|BK006946.2| 322334 - INS 
 tpg|BK006946.2| 766975 + tpg|BK006946.2| 767182 - INS 
 tpg|BK006946.2| 528422 + tpg|BK006946.2| 528311 - INS 
 tpg|BK006946.2| 505103 + tpg|BK006946.2| 505727 - INS 
 tpg|BK006946.2| 638901 + tpg|BK006946.2| 639536 - INS 
 tpg|BK006946.2| 686762 + tpg|BK006946.2| 687121 - INS 
 tpg|BK006946.2| 743932 + tpg|BK006946.2| 743575 - INS 
 tpg|BK006946.2| 753218 + tpg|BK006946.2| 753853 - INS 
 tpg|BK006946.2| 9256 + tpg|BK006946.2| 9866 - INS 
 tpg|BK006946.2| 647382 + tpg|BK006946.2| 647149 - INS 
 tpg|BK006946.2| 182520 + tpg|BK006946.2| 182279 - INS 
 tpg|BK006946.2| 190717 + tpg|BK006946.2| 190577 - INS 
 tpg|BK006946.2| 231531 + tpg|BK006946.2| 232145 - INS 
 tpg|BK006946.2| 897909 + tpg|BK006946.2| 897375 - INS 
 tpg|BK006946.2| 46917 + tpg|BK006946.2| 46494 - INS 
 tpg|BK006946.2| 464161 + tpg|BK006946.2| 463509 - INS 
 tpg|BK006946.2| 463263 + tpg|BK006946.2| 462654 - INS 
 tpg|BK006946.2| 881501 + tpg|BK006946.2| 880903 - INS 
 tpg|BK006946.2| 130651 + tpg|BK006946.2| 130484 - INS 
 tpg|BK006946.2| 431997 + tpg|BK006946.2| 431850 - INS 
 tpg|BK006946.2| 628473 + tpg|BK006946.2| 629107 - INS 
 tpg|BK006946.2| 617730 + tpg|BK006946.2| 618446 - INS 
 tpg|BK006946.2| 426773 + tpg|BK006946.2| 426478 - INS 
 tpg|BK006946.2| 863392 + tpg|BK006946.2| 863840 - INS 
 tpg|BK006946.2| 403708 + tpg|BK006946.2| 403492 - INS 
 tpg|BK006946.2| 640497 + tpg|BK006946.2| 640982 - INS 
 tpg|BK006946.2| 838882 + tpg|BK006946.2| 838792 - INS 
 tpg|BK006946.2| 692368 + tpg|BK006946.2| 692093 - INS 
 tpg|BK006946.2| 814866 + tpg|BK006946.2| 814724 - INS 
 tpg|BK006946.2| 385470 + tpg|BK006946.2| 385065 - INS 
 tpg|BK006946.2| 714256 + tpg|BK006946.2| 714082 - INS 
 tpg|BK006946.2| 713688 + tpg|BK006946.2| 712973 - INS 
 tpg|BK006946.2| 353037 + tpg|BK006946.2| 352690 - INS 
 tpg|BK006946.2| 343655 + tpg|BK006946.2| 343265 - INS 
 tpg|BK006946.2| 103484 + tpg|BK006946.2| 103071 - INS 
 tpg|BK006946.2| 642751 + tpg|BK006946.2| 642725 - INS 
 tpg|BK006946.2| 318408 + tpg|BK006946.2| 318343 - INS 
 tpg|BK006946.2| 837620 + tpg|BK006946.2| 838251 - INS 
 tpg|BK006946.2| 876944 + tpg|BK006946.2| 876672 - INS 
 tpg|BK006946.2| 680540 + tpg|BK006946.2| 680413 - INS 
 tpg|BK006946.2| 647944 + tpg|BK006946.2| 648114 - INS 
 tpg|BK006946.2| 445804 + tpg|BK006946.2| 445892 - INS 
 tpg|BK006946.2| 148825 + tpg|BK006946.2| 149393 - INS 
 tpg|BK006946.2| 671154 + tpg|BK006946.2| 671433 - INS 
 tpg|BK006946.2| 828027 + tpg|BK006946.2| 828584 - INS 
 tpg|BK006946.2| 610589 + tpg|BK006946.2| 610379 - INS 
 tpg|BK006946.2| 153632 + tpg|BK006946.2| 153058 - INS 
 tpg|BK006946.2| 824982 + tpg|BK006946.2| 824909 - INS 
 tpg|BK006946.2| 145876 + tpg|BK006946.2| 145733 - INS 
 tpg|BK006946.2| 919708 + tpg|BK006946.2| 919096 - INS 
 tpg|BK006946.2| 794521 + tpg|BK006946.2| 794514 - INS 
 tpg|BK006946.2| 47795 + tpg|BK006946.2| 48201 - INS 
 tpg|BK006946.2| 302081 + tpg|BK006946.2| 301604 - INS 
 tpg|BK006946.2| 580620 + tpg|BK006946.2| 581346 - INS 
 tpg|BK006946.2| 183452 + tpg|BK006946.2| 182902 - INS 
 tpg|BK006946.2| 339473 + tpg|BK006946.2| 339973 - INS 
 tpg|BK006946.2| 570286 + tpg|BK006946.2| 570783 - INS 
 tpg|BK006946.2| 559440 + tpg|BK006946.2| 559179 - INS 
 tpg|BK006946.2| 751601 + tpg|BK006946.2| 751107 - INS 
 tpg|BK006946.2| 487290 + tpg|BK006946.2| 487942 - INS 
 tpg|BK006946.2| 287026 + tpg|BK006946.2| 286981 - INS 
 tpg|BK006946.2| 922328 + tpg|BK006946.2| 922839 - INS 
 tpg|BK006946.2| 655301 + tpg|BK006946.2| 654799 - INS 
 tpg|BK006946.2| 499078 + tpg|BK006946.2| 498857 - INS 
 tpg|BK006946.2| 776389 + tpg|BK006946.2| 775770 - INS 
 tpg|BK006946.2| 240388 + tpg|BK006946.2| 241022 - INS 
 tpg|BK006946.2| 745934 + tpg|BK006946.2| 746017 - INS 
 tpg|BK006946.2| 446828 + tpg|BK006946.2| 447467 - INS 
 tpg|BK006946.2| 397336 + tpg|BK006946.2| 397981 - INS 
 tpg|BK006946.2| 370638 + tpg|BK006946.2| 371198 - INS 
 tpg|BK006946.2| 332545 + tpg|BK006946.2| 332395 - INS 
 tpg|BK006946.2| 293959 + tpg|BK006946.2| 293860 - INS 
 tpg|BK006946.2| 233828 + tpg|BK006946.2| 233608 - INS 
 tpg|BK006946.2| 599187 + tpg|BK006946.2| 599272 - INS 
 tpg|BK006946.2| 87925 + tpg|BK006946.2| 88510 - INS 
 tpg|BK006946.2| 475645 + tpg|BK006946.2| 475940 - INS 
 tpg|BK006946.2| 28645 + tpg|BK006946.2| 28699 - INS 
 tpg|BK006946.2| 75732 + tpg|BK006946.2| 75200 - INS 
 tpg|BK006946.2| 917045 + tpg|BK006946.2| 916941 - INS 
 tpg|BK006946.2| 323246 + tpg|BK006946.2| 323826 - INS 
 tpg|BK006946.2| 465343 + tpg|BK006946.2| 465271 - INS 
 tpg|BK006946.2| 799775 + tpg|BK006946.2| 800103 - INS 
 tpg|BK006946.2| 689340 + tpg|BK006946.2| 689030 - INS 
 tpg|BK006946.2| 265974 + tpg|BK006946.2| 265877 - INS 
 tpg|BK006946.2| 551772 + tpg|BK006946.2| 551603 - INS 
 tpg|BK006946.2| 184254 + tpg|BK006946.2| 183902 - INS 
 tpg|BK006946.2| 488782 + tpg|BK006946.2| 488554 - INS 
 tpg|BK006946.2| 180002 + tpg|BK006946.2| 180638 - INS 
 tpg|BK006946.2| 310532 + tpg|BK006946.2| 310710 - INS 
 tpg|BK006946.2| 686125 + tpg|BK006946.2| 685695 - INS 
 tpg|BK006946.2| 301291 + tpg|BK006946.2| 300855 - INS 
 tpg|BK006946.2| 510866 + tpg|BK006946.2| 510787 - INS 
 tpg|BK006946.2| 290405 + tpg|BK006946.2| 289747 - INS 
 tpg|BK006946.2| 582612 + tpg|BK006946.2| 582118 - INS 
 tpg|BK006946.2| 682997 + tpg|BK006946.2| 683762 - INS 
 tpg|BK006946.2| 658586 + tpg|BK006946.2| 658392 - INS 
 tpg|BK006946.2| 752309 + tpg|BK006946.2| 751954 - INS 
 tpg|BK006946.2| 810217 + tpg|BK006946.2| 810239 - INS 
 tpg|BK006946.2| 857086 + tpg|BK006946.2| 856717 - INS 
 tpg|BK006946.2| 555507 + tpg|BK006946.2| 555097 - INS 
 tpg|BK006946.2| 893677 + tpg|BK006946.2| 892955 - INS 
 tpg|BK006946.2| 47408 + tpg|BK006946.2| 46910 - INS 
 tpg|BK006946.2| 179467 + tpg|BK006946.2| 179469 - INS 
 tpg|BK006946.2| 144060 + tpg|BK006946.2| 143704 - INS 
 tpg|BK006946.2| 84198 + tpg|BK006946.2| 83990 - INS 
 tpg|BK006946.2| 690872 + tpg|BK006946.2| 690539 - INS 
 tpg|BK006946.2| 891293 + tpg|BK006946.2| 890654 - INS 
 tpg|BK006946.2| 79237 + tpg|BK006946.2| 78883 - INS 
 tpg|BK006946.2| 331196 + tpg|BK006946.2| 330919 - INS 
 tpg|BK006946.2| 630804 + tpg|BK006946.2| 630496 - INS 
 tpg|BK006946.2| 338963 + tpg|BK006946.2| 339290 - INS 
 tpg|BK006946.2| 732052 + tpg|BK006946.2| 731855 - INS 
 tpg|BK006946.2| 49507 + tpg|BK006946.2| 48781 - INS 
 tpg|BK006946.2| 107150 + tpg|BK006946.2| 107151 - INS 
 tpg|BK006946.2| 461787 + tpg|BK006946.2| 461411 - INS 
 tpg|BK006946.2| 210797 + tpg|BK006946.2| 210193 - INS 
 tpg|BK006946.2| 906895 + tpg|BK006946.2| 906789 - INS 
 tpg|BK006946.2| 329923 + tpg|BK006946.2| 329322 - INS 
 tpg|BK006946.2| 252708 + tpg|BK006946.2| 252578 - INS 
 tpg|BK006946.2| 517522 + tpg|BK006946.2| 516853 - INS 
 tpg|BK006946.2| 228364 + tpg|BK006946.2| 228238 - INS 
 tpg|BK006946.2| 365769 + tpg|BK006946.2| 365267 - INS 
 tpg|BK006946.2| 835798 + tpg|BK006946.2| 835700 - INS 
 tpg|BK006946.2| 162165 + tpg|BK006946.2| 161587 - INS 
 tpg|BK006946.2| 596950 + tpg|BK006946.2| 597125 - INS 
 tpg|BK006946.2| 543187 + tpg|BK006946.2| 543195 - INS 
 tpg|BK006946.2| 678604 + tpg|BK006946.2| 678414 - INS 
 tpg|BK006946.2| 56076 + tpg|BK006946.2| 55551 - INS 
 tpg|BK006946.2| 350818 + tpg|BK006946.2| 350379 - INS 
 tpg|BK006946.2| 783823 + tpg|BK006946.2| 783172 - INS 
 tpg|BK006946.2| 89955 + tpg|BK006946.2| 89580 - INS 
 tpg|BK006946.2| 736563 + tpg|BK006946.2| 736503 - INS 
 tpg|BK006946.2| 279355 + tpg|BK006946.2| 279733 - INS 
 tpg|BK006946.2| 563933 + tpg|BK006946.2| 563475 - INS 
 tpg|BK006946.2| 93431 + tpg|BK006946.2| 93008 - INS 
 tpg|BK006946.2| 511666 + tpg|BK006946.2| 511525 - INS 
 tpg|BK006946.2| 91282 + tpg|BK006946.2| 90827 - INS 
 tpg|BK006946.2| 335747 + tpg|BK006946.2| 335201 - INS 
 tpg|BK006946.2| 345737 + tpg|BK006946.2| 345772 - INS 
 tpg|BK006946.2| 698915 + tpg|BK006946.2| 698548 - INS 
 tpg|BK006946.2| 125737 + tpg|BK006946.2| 125682 - INS 
 tpg|BK006946.2| 914605 + tpg|BK006946.2| 914827 - INS 
 tpg|BK006946.2| 132451 + tpg|BK006946.2| 132146 - INS 
 tpg|BK006946.2| 239894 + tpg|BK006946.2| 240579 - INS 
 tpg|BK006946.2| 621654 + tpg|BK006946.2| 621354 - INS 
 tpg|BK006946.2| 497891 + tpg|BK006946.2| 497586 - INS 
 tpg|BK006946.2| 118516 + tpg|BK006946.2| 117876 - INS 
 tpg|BK006946.2| 383172 + tpg|BK006946.2| 382936 - INS 
 tpg|BK006946.2| 256216 + tpg|BK006946.2| 255804 - INS 
 tpg|BK006946.2| 527369 + tpg|BK006946.2| 526806 - INS 
 tpg|BK006946.2| 899134 + tpg|BK006946.2| 899069 - INS 
 tpg|BK006946.2| 733120 + tpg|BK006946.2| 733065 - INS 
 tpg|BK006946.2| 587559 + tpg|BK006946.2| 587168 - INS 
 tpg|BK006946.2| 845387 + tpg|BK006946.2| 844956 - INS 
 tpg|BK006946.2| 480506 + tpg|BK006946.2| 479770 - INS 
 tpg|BK006946.2| 464647 + tpg|BK006946.2| 464455 - INS 
 tpg|BK006946.2| 728306 + tpg|BK006946.2| 727934 - INS 
 tpg|BK006946.2| 139692 + tpg|BK006946.2| 139757 - INS 
 tpg|BK006946.2| 677320 + tpg|BK006946.2| 676694 - INS 
 tpg|BK006946.2| 211787 + tpg|BK006946.2| 211713 - INS 
 tpg|BK006946.2| 502128 + tpg|BK006946.2| 501722 - INS 
 tpg|BK006946.2| 263364 + tpg|BK006946.2| 263449 - INS 
 tpg|BK006946.2| 208227 + tpg|BK006946.2| 207854 - INS 
 tpg|BK006946.2| 91807 + tpg|BK006946.2| 92046 - INS 
 tpg|BK006946.2| 514346 + tpg|BK006946.2| 514297 - INS 
 tpg|BK006946.2| 826324 + tpg|BK006946.2| 825559 - INS 
 tpg|BK006946.2| 366255 + tpg|BK006946.2| 365907 - INS 
 tpg|BK006946.2| 585653 + tpg|BK006946.2| 585646 - INS 
 tpg|BK006946.2| 505609 + tpg|BK006946.2| 506332 - INS 
 tpg|BK006946.2| 602682 + tpg|BK006946.2| 602123 - INS 
 tpg|BK006946.2| 42820 + tpg|BK006946.2| 42511 - INS 
 tpg|BK006946.2| 521224 + tpg|BK006946.2| 520957 - INS 
 tpg|BK006946.2| 883950 + tpg|BK006946.2| 883983 - INS 
 tpg|BK006946.2| 901907 + tpg|BK006946.2| 901946 - INS 
 tpg|BK006946.2| 245909 + tpg|BK006946.2| 245436 - INS 
 tpg|BK006946.2| 877956 + tpg|BK006946.2| 878602 - INS 
 tpg|BK006946.2| 539211 + tpg|BK006946.2| 539465 - INS 
 tpg|BK006946.2| 520120 + tpg|BK006946.2| 519785 - INS 
 tpg|BK006946.2| 709178 + tpg|BK006946.2| 709429 - INS 
 tpg|BK006946.2| 18189 + tpg|BK006946.2| 18192 - INS 
 tpg|BK006946.2| 122454 + tpg|BK006946.2| 122321 - INS 
 tpg|BK006946.2| 734337 + tpg|BK006946.2| 734240 - INS 
 tpg|BK006946.2| 882186 + tpg|BK006946.2| 881509 - INS 
 tpg|BK006946.2| 894104 + tpg|BK006946.2| 893757 - INS 
 tpg|BK006946.2| 27175 + tpg|BK006946.2| 27185 - INS 
 tpg|BK006946.2| 696400 + tpg|BK006946.2| 696143 - INS 
 tpg|BK006946.2| 871409 + tpg|BK006946.2| 872032 - INS 
 tpg|BK006946.2| 333171 + tpg|BK006946.2| 333392 - INS 
 tpg|BK006946.2| 455454 + tpg|BK006946.2| 455297 - INS 
 tpg|BK006946.2| 920870 + tpg|BK006946.2| 920907 - INS 
 tpg|BK006946.2| 437463 + tpg|BK006946.2| 437279 - INS 
 tpg|BK006946.2| 81212 + tpg|BK006946.2| 80843 - INS 
 tpg|BK006946.2| 466470 + tpg|BK006946.2| 465843 - INS 
 tpg|BK006946.2| 243902 + tpg|BK006946.2| 243729 - INS 
 tpg|BK006947.3| 214650 + tpg|BK006947.3| 214674 - INS 
 tpg|BK006947.3| 661500 + tpg|BK006947.3| 661583 - INS 
 tpg|BK006947.3| 226214 + tpg|BK006947.3| 226837 - INS 
 tpg|BK006947.3| 141043 + tpg|BK006947.3| 140679 - INS 
 tpg|BK006947.3| 591086 + tpg|BK006947.3| 590496 - INS 
 tpg|BK006947.3| 528775 + tpg|BK006947.3| 529355 - INS 
 tpg|BK006947.3| 138444 + tpg|BK006947.3| 138732 - INS 
 tpg|BK006947.3| 527891 + tpg|BK006947.3| 528037 - INS 
 tpg|BK006947.3| 210304 + tpg|BK006947.3| 209831 - INS 
 tpg|BK006947.3| 357497 + tpg|BK006947.3| 357025 - INS 
 tpg|BK006947.3| 733965 + tpg|BK006947.3| 733799 - INS 
 tpg|BK006947.3| 298215 + tpg|BK006947.3| 297578 - INS 
 tpg|BK006947.3| 704414 + tpg|BK006947.3| 704478 - INS 
 tpg|BK006947.3| 708050 + tpg|BK006947.3| 707864 - INS 
 tpg|BK006947.3| 455978 + tpg|BK006947.3| 455642 - INS 
 tpg|BK006947.3| 525715 + tpg|BK006947.3| 525298 - INS 
 tpg|BK006947.3| 423186 + tpg|BK006947.3| 423958 - INS 
 tpg|BK006947.3| 540519 + tpg|BK006947.3| 540763 - INS 
 tpg|BK006947.3| 641514 + tpg|BK006947.3| 641221 - INS 
 tpg|BK006947.3| 289616 + tpg|BK006947.3| 289134 - INS 
 tpg|BK006947.3| 702723 + tpg|BK006947.3| 702971 - INS 
 tpg|BK006947.3| 89494 + tpg|BK006947.3| 88899 - INS 
 tpg|BK006947.3| 414031 + tpg|BK006947.3| 413448 - INS T
 tpg|BK006947.3| 465340 + tpg|BK006947.3| 465677 - INS 
 tpg|BK006947.3| 242316 + tpg|BK006947.3| 242016 - INS 
 tpg|BK006947.3| 380214 + tpg|BK006947.3| 379802 - INS 
 tpg|BK006947.3| 506376 + tpg|BK006947.3| 507146 - INS 
 tpg|BK006947.3| 646732 + tpg|BK006947.3| 646487 - INS 
 tpg|BK006947.3| 610272 + tpg|BK006947.3| 610740 - INS 
 tpg|BK006947.3| 207820 + tpg|BK006947.3| 207320 - INS 
 tpg|BK006947.3| 676003 + tpg|BK006947.3| 675430 - INS 
 tpg|BK006947.3| 292877 + tpg|BK006947.3| 293109 - INS 
 tpg|BK006947.3| 630154 + tpg|BK006947.3| 629625 - INS 
 tpg|BK006947.3| 410053 + tpg|BK006947.3| 410012 - INS 
 tpg|BK006947.3| 386059 + tpg|BK006947.3| 386368 - INS 
 tpg|BK006947.3| 757604 + tpg|BK006947.3| 757857 - INS 
 tpg|BK006947.3| 53164 + tpg|BK006947.3| 53325 - INS 
 tpg|BK006947.3| 747091 + tpg|BK006947.3| 747165 - INS 
 tpg|BK006947.3| 440735 + tpg|BK006947.3| 441141 - INS 
 tpg|BK006947.3| 613513 + tpg|BK006947.3| 613449 - INS 
 tpg|BK006947.3| 777254 + tpg|BK006947.3| 777251 - INS 
 tpg|BK006947.3| 534210 + tpg|BK006947.3| 534821 - INS 
 tpg|BK006947.3| 555974 + tpg|BK006947.3| 555940 - INS 
 tpg|BK006947.3| 273318 + tpg|BK006947.3| 272631 - INS 
 tpg|BK006947.3| 686668 + tpg|BK006947.3| 686442 - INS 
 tpg|BK006947.3| 202552 + tpg|BK006947.3| 202652 - INS 
 tpg|BK006947.3| 430065 + tpg|BK006947.3| 430157 - INS 
 tpg|BK006947.3| 332620 + tpg|BK006947.3| 332286 - INS 
 tpg|BK006947.3| 724117 + tpg|BK006947.3| 723590 - INS 
 tpg|BK006947.3| 759409 + tpg|BK006947.3| 758992 - INS 
 tpg|BK006947.3| 674808 + tpg|BK006947.3| 674763 - INS 
 tpg|BK006947.3| 416684 + tpg|BK006947.3| 416246 - INS 
 tpg|BK006947.3| 456809 + tpg|BK006947.3| 456497 - INS 
 tpg|BK006947.3| 480213 + tpg|BK006947.3| 480620 - INS 
 tpg|BK006947.3| 91938 + tpg|BK006947.3| 91826 - INS 
 tpg|BK006936.2| 194812 + tpg|BK006936.2| 195079 - INS 
 tpg|BK006947.3| 684235 + tpg|BK006947.3| 684245 - INS 
 tpg|BK006936.2| 270715 + tpg|BK006936.2| 271014 - INS 
 tpg|BK006947.3| 317628 + tpg|BK006947.3| 317358 - INS 
 tpg|BK006947.3| 311418 + tpg|BK006947.3| 311521 - INS 
 tpg|BK006936.2| 634944 + tpg|BK006936.2| 634832 - INS 
 tpg|BK006947.3| 700601 + tpg|BK006947.3| 700577 - INS 
 tpg|BK006936.2| 106646 + tpg|BK006936.2| 106176 - INS 
 tpg|BK006947.3| 575052 + tpg|BK006947.3| 575324 - INS 
 tpg|BK006947.3| 483675 + tpg|BK006947.3| 483277 - INS 
 tpg|BK006947.3| 492296 + tpg|BK006947.3| 491895 - INS 
 tpg|BK006947.3| 43833 + tpg|BK006947.3| 43137 - INS 
 tpg|BK006936.2| 374003 + tpg|BK006936.2| 373473 - INS 
 tpg|BK006947.3| 479315 + tpg|BK006947.3| 479249 - INS 
 tpg|BK006947.3| 623784 + tpg|BK006947.3| 623948 - INS 
 tpg|BK006936.2| 312316 + tpg|BK006936.2| 311782 - INS 
 tpg|BK006947.3| 643302 + tpg|BK006947.3| 642659 - INS 
 tpg|BK006947.3| 328181 + tpg|BK006947.3| 328397 - INS 
 tpg|BK006947.3| 329629 + tpg|BK006947.3| 329659 - INS 
 tpg|BK006947.3| 690564 + tpg|BK006947.3| 690419 - INS 
 tpg|BK006936.2| 681410 + tpg|BK006936.2| 681711 - INS 
 tpg|BK006947.3| 778541 + tpg|BK006947.3| 779081 - INS 
 tpg|BK006947.3| 337592 + tpg|BK006947.3| 337671 - INS 
 tpg|BK006936.2| 465308 + tpg|BK006936.2| 465222 - INS 
 tpg|BK006947.3| 184190 + tpg|BK006947.3| 183698 - INS 
 tpg|BK006947.3| 502127 + tpg|BK006947.3| 502325 - INS 
 tpg|BK006936.2| 27890 + tpg|BK006936.2| 27627 - INS 
 tpg|BK006947.3| 740365 + tpg|BK006947.3| 740886 - INS 
 tpg|BK006947.3| 195152 + tpg|BK006947.3| 195292 - INS 
 tpg|BK006936.2| 788267 + tpg|BK006936.2| 787770 - INS 
 tpg|BK006936.2| 213099 + tpg|BK006936.2| 212417 - INS 
 tpg|BK006947.3| 315395 + tpg|BK006947.3| 315525 - INS 
 tpg|BK006947.3| 692940 + tpg|BK006947.3| 692956 - INS 
 tpg|BK006947.3| 763108 + tpg|BK006947.3| 763133 - INS 
 tpg|BK006947.3| 780161 + tpg|BK006947.3| 779912 - INS 
 tpg|BK006947.3| 326177 + tpg|BK006947.3| 326843 - INS 
 tpg|BK006947.3| 71354 + tpg|BK006947.3| 70960 - INS 
 tpg|BK006947.3| 265598 + tpg|BK006947.3| 265710 - INS 
 tpg|BK006947.3| 180483 + tpg|BK006947.3| 179754 - INS 
 tpg|BK006936.2| 618761 + tpg|BK006936.2| 619341 - INS 
 tpg|BK006947.3| 189637 + tpg|BK006947.3| 189002 - INS 
 tpg|BK006947.3| 654282 + tpg|BK006947.3| 653820 - INS 
 tpg|BK006947.3| 491064 + tpg|BK006947.3| 490655 - INS 
 tpg|BK006936.2| 244220 + tpg|BK006936.2| 243968 - INS 
 tpg|BK006947.3| 503841 + tpg|BK006947.3| 503091 - INS 
 tpg|BK006947.3| 330191 + tpg|BK006947.3| 330518 - INS 
 tpg|BK006936.2| 176413 + tpg|BK006936.2| 176152 - INS 
 tpg|BK006936.2| 273921 + tpg|BK006936.2| 273634 - INS 
 tpg|BK006947.3| 391264 + tpg|BK006947.3| 391395 - INS 
 tpg|BK006936.2| 247049 + tpg|BK006936.2| 247189 - INS 
 tpg|BK006947.3| 508325 + tpg|BK006947.3| 507804 - INS 
 tpg|BK006936.2| 621796 + tpg|BK006936.2| 621024 - INS 
 tpg|BK006936.2| 117098 + tpg|BK006936.2| 117018 - INS 
 tpg|BK006947.3| 218111 + tpg|BK006947.3| 217905 - INS 
 tpg|BK006936.2| 570299 + tpg|BK006936.2| 570690 - INS 
 tpg|BK006947.3| 363194 + tpg|BK006947.3| 362782 - INS 
 tpg|BK006947.3| 282996 + tpg|BK006947.3| 282559 - INS 
 tpg|BK006947.3| 51618 + tpg|BK006947.3| 51148 - INS 
 tpg|BK006936.2| 314708 + tpg|BK006936.2| 314186 - INS 
 tpg|BK006947.3| 658234 + tpg|BK006947.3| 657689 - INS 
 tpg|BK006936.2| 772062 + tpg|BK006936.2| 771781 - INS 
 tpg|BK006947.3| 216774 + tpg|BK006947.3| 217049 - INS 
 tpg|BK006936.2| 99390 + tpg|BK006936.2| 100008 - INS 
 tpg|BK006936.2| 615699 + tpg|BK006936.2| 615145 - INS 
 tpg|BK006947.3| 701922 + tpg|BK006947.3| 702376 - INS 
 tpg|BK006947.3| 143161 + tpg|BK006947.3| 143353 - INS 
 tpg|BK006936.2| 690781 + tpg|BK006936.2| 690501 - INS 
 tpg|BK006936.2| 761466 + tpg|BK006936.2| 760707 - INS 
 tpg|BK006936.2| 794216 + tpg|BK006936.2| 793841 - INS 
 tpg|BK006947.3| 196149 + tpg|BK006947.3| 196730 - INS 
 tpg|BK006936.2| 422886 + tpg|BK006936.2| 423637 - INS 
 tpg|BK006947.3| 394065 + tpg|BK006947.3| 393953 - INS 
 tpg|BK006947.3| 173180 + tpg|BK006947.3| 173011 - INS 
 tpg|BK006936.2| 649752 + tpg|BK006936.2| 650060 - INS 
 tpg|BK006947.3| 69978 + tpg|BK006947.3| 69852 - INS 
 tpg|BK006947.3| 639675 + tpg|BK006947.3| 639411 - INS 
 tpg|BK006947.3| 756406 + tpg|BK006947.3| 756811 - INS 
 tpg|BK006947.3| 302341 + tpg|BK006947.3| 301935 - INS 
 tpg|BK006947.3| 338193 + tpg|BK006947.3| 338882 - INS 
 tpg|BK006936.2| 193900 + tpg|BK006936.2| 193496 - INS 
 tpg|BK006947.3| 288183 + tpg|BK006947.3| 288296 - INS 
 tpg|BK006947.3| 594412 + tpg|BK006947.3| 594758 - INS 
 tpg|BK006947.3| 120223 + tpg|BK006947.3| 120509 - INS CTATC
 tpg|BK006936.2| 71734 + tpg|BK006936.2| 72457 - INS 
 tpg|BK006947.3| 256595 + tpg|BK006947.3| 256514 - INS 
 tpg|BK006936.2| 526080 + tpg|BK006936.2| 526588 - INS 
 tpg|BK006936.2| 802700 + tpg|BK006936.2| 803414 - INS 
 tpg|BK006947.3| 240823 + tpg|BK006947.3| 240622 - INS 
 tpg|BK006936.2| 237105 + tpg|BK006936.2| 236725 - INS 
 tpg|BK006947.3| 555222 + tpg|BK006947.3| 554673 - INS 
 tpg|BK006936.2| 711952 + tpg|BK006936.2| 711224 - INS 
 tpg|BK006947.3| 547442 + tpg|BK006947.3| 547375 - INS 
 tpg|BK006947.3| 175570 + tpg|BK006947.3| 174991 - INS 
 tpg|BK006936.2| 14049 + tpg|BK006936.2| 13894 - INS 
 tpg|BK006947.3| 37393 + tpg|BK006947.3| 36811 - INS 
 tpg|BK006936.2| 258759 + tpg|BK006936.2| 258833 - INS 
 tpg|BK006947.3| 164335 + tpg|BK006947.3| 165015 - INS 
 tpg|BK006936.2| 518382 + tpg|BK006936.2| 518913 - INS 
 tpg|BK006947.3| 652928 + tpg|BK006947.3| 653230 - INS 
 tpg|BK006947.3| 512765 + tpg|BK006947.3| 512504 - INS 
 tpg|BK006947.3| 736206 + tpg|BK006947.3| 736466 - INS 
 tpg|BK006947.3| 593471 + tpg|BK006947.3| 592952 - INS 
 tpg|BK006947.3| 127847 + tpg|BK006947.3| 127151 - INS 
 tpg|BK006947.3| 392744 + tpg|BK006947.3| 392220 - INS 
 tpg|BK006947.3| 695699 + tpg|BK006947.3| 695400 - INS 
 tpg|BK006947.3| 636876 + tpg|BK006947.3| 637416 - INS 
 tpg|BK006947.3| 286315 + tpg|BK006947.3| 286096 - INS 
 tpg|BK006947.3| 634007 + tpg|BK006947.3| 634559 - INS 
 tpg|BK006947.3| 26286 + tpg|BK006947.3| 25934 - INS 
 tpg|BK006936.2| 433274 + tpg|BK006936.2| 432547 - INS 
 tpg|BK006947.3| 426893 + tpg|BK006947.3| 426824 - INS 
 tpg|BK006947.3| 40533 + tpg|BK006947.3| 40106 - INS 
 tpg|BK006947.3| 59779 + tpg|BK006947.3| 59699 - INS 
 tpg|BK006947.3| 230139 + tpg|BK006947.3| 230709 - INS 
 tpg|BK006947.3| 616825 + tpg|BK006947.3| 616801 - INS 
 tpg|BK006936.2| 19417 + tpg|BK006936.2| 19473 - INS 
 tpg|BK006947.3| 276085 + tpg|BK006947.3| 275822 - INS 
 tpg|BK006936.2| 297303 + tpg|BK006936.2| 297335 - INS 
 tpg|BK006947.3| 343073 + tpg|BK006947.3| 342876 - INS 
 tpg|BK006947.3| 321994 + tpg|BK006947.3| 322522 - INS 
 tpg|BK006936.2| 359371 + tpg|BK006936.2| 359984 - INS 
 tpg|BK006947.3| 205443 + tpg|BK006947.3| 205660 - INS 
 tpg|BK006947.3| 247943 + tpg|BK006947.3| 247308 - INS 
 tpg|BK006947.3| 408538 + tpg|BK006947.3| 408714 - INS 
 tpg|BK006936.2| 133270 + tpg|BK006936.2| 133925 - INS 
 tpg|BK006947.3| 403201 + tpg|BK006947.3| 403483 - INS 
 tpg|BK006936.2| 660406 + tpg|BK006936.2| 661069 - INS 
 tpg|BK006947.3| 531658 + tpg|BK006947.3| 531716 - INS 
 tpg|BK006936.2| 209519 + tpg|BK006936.2| 210287 - INS 
 tpg|BK006947.3| 397778 + tpg|BK006947.3| 398141 - INS 
 tpg|BK006936.2| 593481 + tpg|BK006936.2| 594010 - INS 
 tpg|BK006947.3| 188297 + tpg|BK006947.3| 188164 - INS 
 tpg|BK006936.2| 585470 + tpg|BK006936.2| 584886 - INS 
 tpg|BK006947.3| 371966 + tpg|BK006947.3| 372248 - INS 
 tpg|BK006936.2| 505278 + tpg|BK006936.2| 505551 - INS 
 tpg|BK006947.3| 509071 + tpg|BK006947.3| 508784 - INS 
 tpg|BK006947.3| 667806 + tpg|BK006947.3| 668370 - INS 
 tpg|BK006947.3| 476648 + tpg|BK006947.3| 476170 - INS 
 tpg|BK006936.2| 529649 + tpg|BK006936.2| 529612 - INS 
 tpg|BK006947.3| 212573 + tpg|BK006947.3| 212626 - INS 
 tpg|BK006945.2| 1031456 + tpg|BK006945.2| 1031958 - INS 
 tpg|BK006936.2| 445209 + tpg|BK006936.2| 444876 - INS 
 tpg|BK006947.3| 541817 + tpg|BK006947.3| 541983 - INS 
 tpg|BK006936.2| 370204 + tpg|BK006936.2| 370173 - INS 
 tpg|BK006936.2| 302904 + tpg|BK006936.2| 302280 - INS 
 tpg|BK006947.3| 543252 + tpg|BK006947.3| 543236 - INS 
 tpg|BK006936.2| 316712 + tpg|BK006936.2| 317306 - INS 
 tpg|BK006947.3| 697889 + tpg|BK006947.3| 697370 - INS 
 tpg|BK006945.2| 97797 + tpg|BK006945.2| 97971 - INS 
 tpg|BK006936.2| 773688 + tpg|BK006936.2| 774222 - INS 
 tpg|BK006947.3| 781182 + tpg|BK006947.3| 781331 - INS 
 tpg|BK006947.3| 161179 + tpg|BK006947.3| 160521 - INS 
 tpg|BK006936.2| 59893 + tpg|BK006936.2| 59504 - INS 
 tpg|BK006945.2| 165169 + tpg|BK006945.2| 165726 - INS 
 tpg|BK006947.3| 160159 + tpg|BK006947.3| 159683 - INS 
 tpg|BK006936.2| 687131 + tpg|BK006936.2| 687286 - INS 
 tpg|BK006947.3| 727727 + tpg|BK006947.3| 727378 - INS 
 tpg|BK006945.2| 237660 + tpg|BK006945.2| 236908 - INS 
 tpg|BK006936.2| 629369 + tpg|BK006936.2| 629229 - INS 
 tpg|BK006947.3| 65474 + tpg|BK006947.3| 65434 - INS 
 tpg|BK006947.3| 349934 + tpg|BK006947.3| 349547 - INS 
 tpg|BK006947.3| 354521 + tpg|BK006947.3| 354729 - INS 
 tpg|BK006936.2| 755326 + tpg|BK006936.2| 754855 - INS 
 tpg|BK006945.2| 560064 + tpg|BK006945.2| 560792 - INS 
 tpg|BK006947.3| 145401 + tpg|BK006947.3| 145706 - INS 
 tpg|BK006947.3| 85630 + tpg|BK006947.3| 86367 - INS 
 tpg|BK006947.3| 375324 + tpg|BK006947.3| 374974 - INS 
 tpg|BK006936.2| 164268 + tpg|BK006936.2| 165040 - INS 
 tpg|BK006945.2| 36685 + tpg|BK006945.2| 36599 - INS 
 tpg|BK006947.3| 680533 + tpg|BK006947.3| 680789 - INS 
 tpg|BK006947.3| 721046 + tpg|BK006947.3| 720551 - INS 
 tpg|BK006947.3| 581670 + tpg|BK006947.3| 582292 - INS 
 tpg|BK006945.2| 388721 + tpg|BK006945.2| 389323 - INS 
 tpg|BK006947.3| 73611 + tpg|BK006947.3| 74296 - INS 
 tpg|BK006947.3| 63578 + tpg|BK006947.3| 63323 - INS 
 tpg|BK006947.3| 93428 + tpg|BK006947.3| 92861 - INS 
 tpg|BK006945.2| 280407 + tpg|BK006945.2| 280063 - INS 
 tpg|BK006947.3| 31045 + tpg|BK006947.3| 30809 - INS 
 tpg|BK006947.3| 80776 + tpg|BK006947.3| 81177 - INS 
 tpg|BK006945.2| 326292 + tpg|BK006945.2| 326708 - INS 
 tpg|BK006936.2| 24621 + tpg|BK006936.2| 24852 - INS 
 tpg|BK006945.2| 512696 + tpg|BK006945.2| 512599 - INS 
 tpg|BK006945.2| 923215 + tpg|BK006945.2| 923010 - INS 
 tpg|BK006947.3| 94421 + tpg|BK006947.3| 93871 - INS 
 tpg|BK006945.2| 260828 + tpg|BK006945.2| 260521 - INS 
 tpg|BK006947.3| 443975 + tpg|BK006947.3| 443950 - INS 
 tpg|BK006945.2| 962670 + tpg|BK006945.2| 962617 - INS 
 tpg|BK006936.2| 531300 + tpg|BK006936.2| 531593 - INS 
 tpg|BK006947.3| 95966 + tpg|BK006947.3| 95722 - INS 
 tpg|BK006936.2| 709920 + tpg|BK006936.2| 709764 - INS 
 tpg|BK006947.3| 42279 + tpg|BK006947.3| 42113 - INS 
 tpg|BK006945.2| 661890 + tpg|BK006945.2| 662320 - INS 
 tpg|BK006947.3| 45161 + tpg|BK006947.3| 45705 - INS 
 tpg|BK006936.2| 630471 + tpg|BK006936.2| 631003 - INS 
 tpg|BK006945.2| 553652 + tpg|BK006945.2| 553396 - INS 
 tpg|BK006936.2| 49343 + tpg|BK006936.2| 49792 - INS 
 tpg|BK006947.3| 660596 + tpg|BK006947.3| 660298 - INS 
 tpg|BK006947.3| 385320 + tpg|BK006947.3| 384589 - INS 
 tpg|BK006936.2| 777643 + tpg|BK006936.2| 777058 - INS 
 tpg|BK006945.2| 558302 + tpg|BK006945.2| 559052 - INS 
 tpg|BK006947.3| 105054 + tpg|BK006947.3| 104885 - INS 
 tpg|BK006936.2| 341208 + tpg|BK006936.2| 341520 - INS 
 tpg|BK006947.3| 720091 + tpg|BK006947.3| 719591 - INS 
 tpg|BK006936.2| 350061 + tpg|BK006936.2| 349912 - INS 
 tpg|BK006945.2| 514320 + tpg|BK006945.2| 513975 - INS 
 tpg|BK006947.3| 719527 + tpg|BK006947.3| 719021 - INS 
 tpg|BK006936.2| 204128 + tpg|BK006936.2| 204035 - INS 
 tpg|BK006947.3| 650259 + tpg|BK006947.3| 649815 - INS 
 tpg|BK006945.2| 1017707 + tpg|BK006945.2| 1018215 - INS 
 tpg|BK006936.2| 364659 + tpg|BK006936.2| 364745 - INS 
 tpg|BK006947.3| 458294 + tpg|BK006947.3| 458256 - INS 
 tpg|BK006947.3| 648941 + tpg|BK006947.3| 648841 - INS 
 tpg|BK006936.2| 494840 + tpg|BK006936.2| 494987 - INS 
 tpg|BK006947.3| 691933 + tpg|BK006947.3| 691373 - INS 
 tpg|BK006947.3| 431086 + tpg|BK006947.3| 431847 - INS 
 tpg|BK006947.3| 106474 + tpg|BK006947.3| 105998 - INS 
 tpg|BK006945.2| 969239 + tpg|BK006945.2| 969782 - INS 
 tpg|BK006947.3| 651399 + tpg|BK006947.3| 651077 - INS 
 tpg|BK006945.2| 735414 + tpg|BK006945.2| 735434 - INS 
 tpg|BK006947.3| 770268 + tpg|BK006947.3| 770759 - INS 
 tpg|BK006936.2| 390320 + tpg|BK006936.2| 390861 - INS 
 tpg|BK006945.2| 757378 + tpg|BK006945.2| 757989 - INS 
 tpg|BK006936.2| 162318 + tpg|BK006936.2| 161645 - INS 
 tpg|BK006947.3| 314444 + tpg|BK006947.3| 314024 - INS 
 tpg|BK006936.2| 146542 + tpg|BK006936.2| 145985 - INS 
 tpg|BK006947.3| 290349 + tpg|BK006947.3| 290492 - INS 
 tpg|BK006945.2| 281954 + tpg|BK006945.2| 282507 - INS 
 tpg|BK006947.3| 21317 + tpg|BK006947.3| 21388 - INS 
 tpg|BK006936.2| 45477 + tpg|BK006936.2| 45219 - INS 
 tpg|BK006945.2| 367562 + tpg|BK006945.2| 368046 - INS 
 tpg|BK006947.3| 87640 + tpg|BK006947.3| 87104 - INS 
 tpg|BK006947.3| 609100 + tpg|BK006947.3| 608721 - INS 
 tpg|BK006936.2| 299499 + tpg|BK006936.2| 299393 - INS 
 tpg|BK006947.3| 679760 + tpg|BK006947.3| 679485 - INS 
 tpg|BK006936.2| 544903 + tpg|BK006936.2| 544423 - INS 
 tpg|BK006945.2| 385869 + tpg|BK006945.2| 385720 - INS 
 tpg|BK006947.3| 618994 + tpg|BK006947.3| 618878 - INS 
 tpg|BK006947.3| 299514 + tpg|BK006947.3| 299084 - INS 
 tpg|BK006936.2| 313345 + tpg|BK006936.2| 313136 - INS 
 tpg|BK006945.2| 970685 + tpg|BK006945.2| 970505 - INS 
 tpg|BK006947.3| 454357 + tpg|BK006947.3| 454513 - INS 
 tpg|BK006947.3| 533588 + tpg|BK006947.3| 533499 - INS 
 tpg|BK006945.2| 340960 + tpg|BK006945.2| 341712 - INS 
 tpg|BK006947.3| 633418 + tpg|BK006947.3| 632685 - INS 
 tpg|BK006936.2| 379554 + tpg|BK006936.2| 379120 - INS 
 tpg|BK006945.2| 958811 + tpg|BK006945.2| 959575 - INS 
 tpg|BK006947.3| 708922 + tpg|BK006947.3| 708861 - INS 
 tpg|BK006936.2| 434134 + tpg|BK006936.2| 434306 - INS 
 tpg|BK006936.2| 706725 + tpg|BK006936.2| 707173 - INS 
 tpg|BK006945.2| 191795 + tpg|BK006945.2| 192104 - INS 
 tpg|BK006936.2| 692640 + tpg|BK006936.2| 693109 - INS 
 tpg|BK006936.2| 231137 + tpg|BK006936.2| 230369 - INS 
 tpg|BK006945.2| 281357 + tpg|BK006945.2| 280849 - INS 
 tpg|BK006936.2| 601246 + tpg|BK006936.2| 601891 - INS 
 tpg|BK006947.3| 743169 + tpg|BK006947.3| 743622 - INS 
 tpg|BK006945.2| 575005 + tpg|BK006945.2| 574429 - INS 
 tpg|BK006936.2| 527569 + tpg|BK006936.2| 527807 - INS 
 tpg|BK006947.3| 49652 + tpg|BK006947.3| 50165 - INS 
 tpg|BK006947.3| 156920 + tpg|BK006947.3| 156868 - INS 
 tpg|BK006936.2| 315431 + tpg|BK006936.2| 315421 - INS AA
 tpg|BK006947.3| 738130 + tpg|BK006947.3| 737654 - INS 
 tpg|BK006947.3| 461315 + tpg|BK006947.3| 461127 - INS 
 tpg|BK006936.2| 309806 + tpg|BK006936.2| 309317 - INS 
 tpg|BK006945.2| 94677 + tpg|BK006945.2| 94663 - INS 
 tpg|BK006947.3| 517178 + tpg|BK006947.3| 517812 - INS 
 tpg|BK006947.3| 38195 + tpg|BK006947.3| 38532 - INS 
 tpg|BK006936.2| 332990 + tpg|BK006936.2| 333147 - INS 
 tpg|BK006947.3| 450220 + tpg|BK006947.3| 449978 - INS 
 tpg|BK006945.2| 288232 + tpg|BK006945.2| 288624 - INS 
 tpg|BK006947.3| 228259 + tpg|BK006947.3| 228799 - INS 
 tpg|BK006947.3| 518656 + tpg|BK006947.3| 518519 - INS 
 tpg|BK006947.3| 728981 + tpg|BK006947.3| 728956 - INS 
 tpg|BK006947.3| 57477 + tpg|BK006947.3| 57130 - INS 
 tpg|BK006945.2| 195501 + tpg|BK006945.2| 195550 - INS 
 tpg|BK006947.3| 550084 + tpg|BK006947.3| 550088 - INS 
 tpg|BK006947.3| 243841 + tpg|BK006947.3| 244084 - INS 
 tpg|BK006945.2| 291135 + tpg|BK006945.2| 290962 - INS 
 tpg|BK006947.3| 204202 + tpg|BK006947.3| 203756 - INS 
 tpg|BK006945.2| 78788 + tpg|BK006945.2| 78450 - INS 
 tpg|BK006947.3| 585493 + tpg|BK006947.3| 585291 - INS 
 tpg|BK006936.2| 207058 + tpg|BK006936.2| 207169 - INS TT
 tpg|BK006947.3| 152339 + tpg|BK006947.3| 152972 - INS 
 tpg|BK006945.2| 625813 + tpg|BK006945.2| 625550 - INS 
 tpg|BK006947.3| 389194 + tpg|BK006947.3| 389472 - INS 
 tpg|BK006947.3| 679069 + tpg|BK006947.3| 678933 - INS 
 tpg|BK006945.2| 752004 + tpg|BK006945.2| 751285 - INS 
 tpg|BK006936.2| 685825 + tpg|BK006936.2| 686018 - INS 
 tpg|BK006947.3| 267262 + tpg|BK006947.3| 267552 - INS 
 tpg|BK006945.2| 204320 + tpg|BK006945.2| 203608 - INS 
 tpg|BK006947.3| 751964 + tpg|BK006947.3| 752448 - INS 
 tpg|BK006936.2| 65570 + tpg|BK006936.2| 65607 - INS 
 tpg|BK006947.3| 172411 + tpg|BK006947.3| 172338 - INS 
 tpg|BK006945.2| 30454 + tpg|BK006945.2| 30071 - INS 
 tpg|BK006947.3| 358788 + tpg|BK006947.3| 358729 - INS 
 tpg|BK006936.2| 199009 + tpg|BK006936.2| 198790 - INS 
 tpg|BK006945.2| 366180 + tpg|BK006945.2| 366217 - INS 
 tpg|BK006947.3| 350463 + tpg|BK006947.3| 351102 - INS 
 tpg|BK006936.2| 571678 + tpg|BK006936.2| 572308 - INS 
 tpg|BK006936.2| 87302 + tpg|BK006936.2| 86689 - INS 
 tpg|BK006945.2| 391613 + tpg|BK006945.2| 391831 - INS 
 tpg|BK006947.3| 291646 + tpg|BK006947.3| 292136 - INS 
 tpg|BK006947.3| 614273 + tpg|BK006947.3| 614439 - INS 
 tpg|BK006945.2| 169522 + tpg|BK006945.2| 169296 - INS 
 tpg|BK006936.2| 393984 + tpg|BK006936.2| 394253 - INS 
 tpg|BK006947.3| 296506 + tpg|BK006947.3| 295779 - INS 
 tpg|BK006945.2| 418745 + tpg|BK006945.2| 418800 - INS 
 tpg|BK006947.3| 333954 + tpg|BK006947.3| 334228 - INS 
 tpg|BK006936.2| 367654 + tpg|BK006936.2| 367065 - INS 
 tpg|BK006947.3| 321065 + tpg|BK006947.3| 320774 - INS 
 tpg|BK006945.2| 103620 + tpg|BK006945.2| 103185 - INS 
 tpg|BK006947.3| 306189 + tpg|BK006947.3| 305519 - INS 
 tpg|BK006947.3| 630841 + tpg|BK006947.3| 631447 - INS 
 tpg|BK006936.2| 372791 + tpg|BK006936.2| 372034 - INS 
 tpg|BK006945.2| 23892 + tpg|BK006945.2| 24201 - INS 
 tpg|BK006947.3| 742381 + tpg|BK006947.3| 742322 - INS 
 tpg|BK006947.3| 184890 + tpg|BK006947.3| 184588 - INS 
 tpg|BK006936.2| 236275 + tpg|BK006936.2| 235881 - INS 
 tpg|BK006947.3| 401525 + tpg|BK006947.3| 401460 - INS 
 tpg|BK006947.3| 527161 + tpg|BK006947.3| 526867 - INS 
 tpg|BK006936.2| 107546 + tpg|BK006936.2| 107003 - INS 
 tpg|BK006945.2| 382681 + tpg|BK006945.2| 382456 - INS 
 tpg|BK006947.3| 224687 + tpg|BK006947.3| 224431 - INS 
 tpg|BK006936.2| 94509 + tpg|BK006936.2| 95252 - INS 
 tpg|BK006947.3| 422326 + tpg|BK006947.3| 422767 - INS 
 tpg|BK006945.2| 346913 + tpg|BK006945.2| 346800 - INS 
 tpg|BK006947.3| 435282 + tpg|BK006947.3| 434939 - INS 
 tpg|BK006936.2| 451432 + tpg|BK006936.2| 451435 - INS 
 tpg|BK006947.3| 125744 + tpg|BK006947.3| 125652 - INS 
 tpg|BK006947.3| 132533 + tpg|BK006947.3| 132189 - INS 
 tpg|BK006936.2| 624176 + tpg|BK006936.2| 623484 - INS 
 tpg|BK006947.3| 133887 + tpg|BK006947.3| 134586 - INS 
 tpg|BK006936.2| 583900 + tpg|BK006936.2| 583467 - INS 
 tpg|BK006947.3| 635746 + tpg|BK006947.3| 636486 - INS 
 tpg|BK006947.3| 725063 + tpg|BK006947.3| 725442 - INS 
 tpg|BK006945.2| 617761 + tpg|BK006945.2| 617128 - INS 
 tpg|BK006936.2| 749619 + tpg|BK006936.2| 749462 - INS 
 tpg|BK006947.3| 762291 + tpg|BK006947.3| 761684 - INS 
 tpg|BK006945.2| 325516 + tpg|BK006945.2| 325185 - INS 
 tpg|BK006936.2| 414642 + tpg|BK006936.2| 414413 - INS 
 tpg|BK006947.3| 761208 + tpg|BK006947.3| 761144 - INS 
 tpg|BK006945.2| 893557 + tpg|BK006945.2| 893397 - INS 
 tpg|BK006947.3| 34423 + tpg|BK006947.3| 33846 - INS 
 tpg|BK006936.2| 750352 + tpg|BK006936.2| 750932 - INS 
 tpg|BK006947.3| 322961 + tpg|BK006947.3| 322989 - INS 
 tpg|BK006947.3| 439474 + tpg|BK006947.3| 440161 - INS 
 tpg|BK006947.3| 767293 + tpg|BK006947.3| 766764 - INS 
 tpg|BK006947.3| 166944 + tpg|BK006947.3| 167128 - INS 
 tpg|BK006945.2| 370433 + tpg|BK006945.2| 369958 - INS 
 tpg|BK006947.3| 671069 + tpg|BK006947.3| 670636 - INS 
 tpg|BK006945.2| 783890 + tpg|BK006945.2| 783411 - INS 
 tpg|BK006947.3| 666150 + tpg|BK006947.3| 665947 - INS 
 tpg|BK006945.2| 716188 + tpg|BK006945.2| 716568 - INS 
 tpg|BK006947.3| 746129 + tpg|BK006947.3| 746574 - INS 
 tpg|BK006947.3| 124544 + tpg|BK006947.3| 124097 - INS 
 tpg|BK006945.2| 327527 + tpg|BK006945.2| 327498 - INS 
 tpg|BK006947.3| 115958 + tpg|BK006947.3| 115869 - INS 
 tpg|BK006947.3| 129425 + tpg|BK006947.3| 128895 - INS 
 tpg|BK006947.3| 114993 + tpg|BK006947.3| 114680 - INS 
 tpg|BK006945.2| 50069 + tpg|BK006945.2| 49435 - INS 
 tpg|BK006947.3| 580369 + tpg|BK006947.3| 580903 - INS 
 tpg|BK006947.3| 81368 + tpg|BK006947.3| 81577 - INS 
 tpg|BK006945.2| 1064858 + tpg|BK006945.2| 1064442 - INS 
 tpg|BK006947.3| 373450 + tpg|BK006947.3| 372806 - INS 
 tpg|BK006947.3| 706318 + tpg|BK006947.3| 706937 - INS 
 tpg|BK006947.3| 441968 + tpg|BK006947.3| 441926 - INS 
 tpg|BK006947.3| 735581 + tpg|BK006947.3| 735021 - INS 
 tpg|BK006945.2| 705363 + tpg|BK006945.2| 704848 - INS 
 tpg|BK006947.3| 374385 + tpg|BK006947.3| 373614 - INS 
 tpg|BK006945.2| 424074 + tpg|BK006945.2| 423963 - INS 
 tpg|BK006947.3| 516632 + tpg|BK006947.3| 515992 - INS 
 tpg|BK006945.2| 792634 + tpg|BK006945.2| 792064 - INS 
 tpg|BK006947.3| 772632 + tpg|BK006947.3| 771982 - INS 
 tpg|BK006947.3| 364972 + tpg|BK006947.3| 364436 - INS 
 tpg|BK006945.2| 682582 + tpg|BK006945.2| 682117 - INS 
 tpg|BK006947.3| 407195 + tpg|BK006947.3| 406734 - INS 
 tpg|BK006947.3| 201821 + tpg|BK006947.3| 201359 - INS 
 tpg|BK006947.3| 109347 + tpg|BK006947.3| 109129 - INS 
 tpg|BK006945.2| 903666 + tpg|BK006945.2| 904078 - INS 
 tpg|BK006947.3| 470279 + tpg|BK006947.3| 469920 - INS 
 tpg|BK006947.3| 669807 + tpg|BK006947.3| 669191 - INS 
 tpg|BK006945.2| 354464 + tpg|BK006945.2| 354658 - INS 
 tpg|BK006947.3| 395403 + tpg|BK006947.3| 395060 - INS 
 tpg|BK006945.2| 72663 + tpg|BK006945.2| 72746 - INS 
 tpg|BK006945.2| 279047 + tpg|BK006945.2| 279688 - INS 
 tpg|BK006936.2| 266458 + tpg|BK006936.2| 265962 - INS 
 tpg|BK006945.2| 338195 + tpg|BK006945.2| 337769 - INS 
 tpg|BK006945.2| 501252 + tpg|BK006945.2| 501582 - INS 
 tpg|BK006947.3| 464316 + tpg|BK006947.3| 463569 - INS 
 tpg|BK006936.2| 409127 + tpg|BK006936.2| 408492 - INS 
 tpg|BK006945.2| 887243 + tpg|BK006945.2| 888015 - INS 
 tpg|BK006936.2| 680082 + tpg|BK006936.2| 679336 - INS 
 tpg|BK006947.3| 91011 + tpg|BK006947.3| 91139 - INS 
 tpg|BK006936.2| 77038 + tpg|BK006936.2| 76484 - INS 
 tpg|BK006947.3| 404285 + tpg|BK006947.3| 404096 - INS 
 tpg|BK006947.3| 457461 + tpg|BK006947.3| 457147 - INS 
 tpg|BK006947.3| 215626 + tpg|BK006947.3| 216309 - INS 
 tpg|BK006945.2| 399634 + tpg|BK006945.2| 399696 - INS 
 tpg|BK006947.3| 689405 + tpg|BK006947.3| 688934 - INS 
 tpg|BK006947.3| 219550 + tpg|BK006947.3| 219735 - INS 
 tpg|BK006945.2| 403217 + tpg|BK006945.2| 403149 - INS 
 tpg|BK006947.3| 672327 + tpg|BK006947.3| 672308 - INS 
 tpg|BK006945.2| 422219 + tpg|BK006945.2| 422288 - INS 
 tpg|BK006936.2| 509722 + tpg|BK006936.2| 508981 - INS 
 tpg|BK006947.3| 750085 + tpg|BK006947.3| 750380 - INS 
 tpg|BK006947.3| 452912 + tpg|BK006947.3| 453275 - INS 
 tpg|BK006936.2| 790335 + tpg|BK006936.2| 790490 - INS 
 tpg|BK006947.3| 444994 + tpg|BK006947.3| 444977 - INS 
 tpg|BK006936.2| 167304 + tpg|BK006936.2| 166835 - INS 
 tpg|BK006945.2| 54393 + tpg|BK006945.2| 54339 - INS 
 tpg|BK006936.2| 140065 + tpg|BK006936.2| 139312 - INS 
 tpg|BK006945.2| 498367 + tpg|BK006945.2| 498891 - INS 
 tpg|BK006947.3| 752750 + tpg|BK006947.3| 752917 - INS 
 tpg|BK006936.2| 130899 + tpg|BK006936.2| 130581 - INS 
 tpg|BK006947.3| 168333 + tpg|BK006947.3| 168373 - INS 
 tpg|BK006945.2| 361123 + tpg|BK006945.2| 360605 - INS 
 tpg|BK006936.2| 550691 + tpg|BK006936.2| 550532 - INS 
 tpg|BK006936.2| 492714 + tpg|BK006936.2| 492943 - INS 
 tpg|BK006945.2| 963462 + tpg|BK006945.2| 963536 - INS 
 tpg|BK006947.3| 748017 + tpg|BK006947.3| 747968 - INS 
 tpg|BK006936.2| 86050 + tpg|BK006936.2| 85543 - INS 
 tpg|BK006947.3| 76262 + tpg|BK006947.3| 76633 - INS 
 tpg|BK006945.2| 534353 + tpg|BK006945.2| 534199 - INS 
 tpg|BK006936.2| 419558 + tpg|BK006936.2| 419295 - INS 
 tpg|BK006947.3| 32163 + tpg|BK006947.3| 31539 - INS 
 tpg|BK006945.2| 826167 + tpg|BK006945.2| 825533 - INS 
 tpg|BK006947.3| 148352 + tpg|BK006947.3| 148289 - INS 
 tpg|BK006947.3| 274098 + tpg|BK006947.3| 273658 - INS 
 tpg|BK006936.2| 203143 + tpg|BK006936.2| 203448 - INS 
 tpg|BK006947.3| 345928 + tpg|BK006947.3| 346223 - INS 
 tpg|BK006947.3| 72462 + tpg|BK006947.3| 72702 - INS 
 tpg|BK006947.3| 19123 + tpg|BK006947.3| 19712 - INS 
 tpg|BK006936.2| 659417 + tpg|BK006936.2| 659264 - INS 
 tpg|BK006947.3| 710452 + tpg|BK006947.3| 710858 - INS 
 tpg|BK006936.2| 557437 + tpg|BK006936.2| 557130 - INS 
 tpg|BK006947.3| 131821 + tpg|BK006947.3| 131379 - INS 
 tpg|BK006945.2| 267081 + tpg|BK006945.2| 267543 - INS 
 tpg|BK006936.2| 336542 + tpg|BK006936.2| 336619 - INS 
 tpg|BK006947.3| 82537 + tpg|BK006947.3| 82961 - INS 
 tpg|BK006947.3| 306934 + tpg|BK006947.3| 306444 - INS 
 tpg|BK006936.2| 654524 + tpg|BK006936.2| 653949 - INS 
 tpg|BK006945.2| 838798 + tpg|BK006945.2| 839357 - INS 
 tpg|BK006936.2| 205711 + tpg|BK006936.2| 206222 - INS 
 tpg|BK006947.3| 560535 + tpg|BK006947.3| 560096 - INS 
 tpg|BK006936.2| 721199 + tpg|BK006936.2| 720641 - INS 
 tpg|BK006947.3| 551262 + tpg|BK006947.3| 550918 - INS 
 tpg|BK006945.2| 157280 + tpg|BK006945.2| 156799 - INS 
 tpg|BK006947.3| 619943 + tpg|BK006947.3| 619820 - INS 
 tpg|BK006947.3| 169544 + tpg|BK006947.3| 170111 - INS 
 tpg|BK006947.3| 295253 + tpg|BK006947.3| 294719 - INS 
 tpg|BK006936.2| 481766 + tpg|BK006936.2| 481299 - INS 
 tpg|BK006947.3| 282314 + tpg|BK006947.3| 281820 - INS 
 tpg|BK006936.2| 691889 + tpg|BK006936.2| 691741 - INS 
 tpg|BK006947.3| 183053 + tpg|BK006947.3| 182584 - INS 
 tpg|BK006945.2| 715127 + tpg|BK006945.2| 715014 - INS 
 tpg|BK006936.2| 459687 + tpg|BK006936.2| 459876 - INS 
 tpg|BK006947.3| 497418 + tpg|BK006947.3| 497575 - INS 
 tpg|BK006947.3| 498954 + tpg|BK006947.3| 498209 - INS 
 tpg|BK006945.2| 649262 + tpg|BK006945.2| 648721 - INS 
 tpg|BK006947.3| 270543 + tpg|BK006947.3| 270335 - INS 
 tpg|BK006936.2| 701325 + tpg|BK006936.2| 701503 - INS 
 tpg|BK006947.3| 68895 + tpg|BK006947.3| 68999 - INS 
 tpg|BK006936.2| 252880 + tpg|BK006936.2| 253219 - INS 
 tpg|BK006945.2| 849739 + tpg|BK006945.2| 849591 - INS 
 tpg|BK006945.2| 161550 + tpg|BK006945.2| 160983 - INS 
 tpg|BK006947.3| 687666 + tpg|BK006947.3| 687249 - INS 
 tpg|BK006947.3| 625919 + tpg|BK006947.3| 625780 - INS 
 tpg|BK006945.2| 712995 + tpg|BK006945.2| 713312 - INS 
 tpg|BK006947.3| 383065 + tpg|BK006947.3| 383803 - INS 
 tpg|BK006936.2| 267332 + tpg|BK006936.2| 267614 - INS 
 tpg|BK006947.3| 730277 + tpg|BK006947.3| 730670 - INS 
 tpg|BK006936.2| 564183 + tpg|BK006936.2| 563933 - INS 
 tpg|BK006945.2| 151876 + tpg|BK006945.2| 152439 - INS 
 tpg|BK006947.3| 271709 + tpg|BK006947.3| 271619 - INS 
 tpg|BK006936.2| 447777 + tpg|BK006936.2| 448144 - INS 
 tpg|BK006947.3| 381607 + tpg|BK006947.3| 380990 - INS 
 tpg|BK006947.3| 303705 + tpg|BK006947.3| 304077 - INS 
 tpg|BK006945.2| 628739 + tpg|BK006945.2| 628401 - INS 
 tpg|BK006936.2| 684497 + tpg|BK006936.2| 684768 - INS 
 tpg|BK006947.3| 387560 + tpg|BK006947.3| 387387 - INS 
 tpg|BK006947.3| 28129 + tpg|BK006947.3| 27376 - INS 
 tpg|BK006936.2| 149032 + tpg|BK006936.2| 149745 - INS 
 tpg|BK006947.3| 557158 + tpg|BK006947.3| 556642 - INS 
 tpg|BK006945.2| 351963 + tpg|BK006945.2| 351401 - INS 
 tpg|BK006945.2| 841586 + tpg|BK006945.2| 841690 - INS 
 tpg|BK006936.2| 439819 + tpg|BK006936.2| 439422 - INS 
 tpg|BK006947.3| 583147 + tpg|BK006947.3| 582915 - INS 
 tpg|BK006947.3| 35317 + tpg|BK006947.3| 35482 - INS 
 tpg|BK006936.2| 457031 + tpg|BK006936.2| 457084 - INS 
 tpg|BK006945.2| 729012 + tpg|BK006945.2| 729551 - INS 
 tpg|BK006947.3| 56123 + tpg|BK006947.3| 56374 - INS 
 tpg|BK006947.3| 232268 + tpg|BK006947.3| 231686 - INS 
 tpg|BK006945.2| 863510 + tpg|BK006945.2| 862777 - INS 
 tpg|BK006947.3| 29058 + tpg|BK006947.3| 28895 - INS 
 tpg|BK006947.3| 448796 + tpg|BK006947.3| 448167 - INS 
 tpg|BK006947.3| 459730 + tpg|BK006947.3| 459453 - INS AAAGA
 tpg|BK006945.2| 853523 + tpg|BK006945.2| 853555 - INS 
 tpg|BK006936.2| 56753 + tpg|BK006936.2| 56378 - INS 
 tpg|BK006936.2| 762266 + tpg|BK006936.2| 761697 - INS 
 tpg|BK006947.3| 776310 + tpg|BK006947.3| 776017 - INS 
 tpg|BK006947.3| 261949 + tpg|BK006947.3| 262325 - INS 
 tpg|BK006947.3| 716595 + tpg|BK006947.3| 716742 - INS 
 tpg|BK006947.3| 715081 + tpg|BK006947.3| 714908 - INS 
 tpg|BK006947.3| 225217 + tpg|BK006947.3| 225127 - INS 
 tpg|BK006936.2| 735639 + tpg|BK006936.2| 736154 - INS 
 tpg|BK006947.3| 252231 + tpg|BK006947.3| 251879 - INS 
 tpg|BK006945.2| 81702 + tpg|BK006945.2| 81409 - INS 
 tpg|BK006947.3| 84890 + tpg|BK006947.3| 85622 - INS 
 tpg|BK006936.2| 160224 + tpg|BK006936.2| 160478 - INS 
 tpg|BK006947.3| 242930 + tpg|BK006947.3| 242787 - INS 
 tpg|BK006936.2| 573780 + tpg|BK006936.2| 573805 - INS 
 tpg|BK006947.3| 433483 + tpg|BK006947.3| 433082 - INS 
 tpg|BK006936.2| 35865 + tpg|BK006936.2| 36155 - INS 
 tpg|BK006947.3| 163585 + tpg|BK006947.3| 163968 - INS 
 tpg|BK006936.2| 513873 + tpg|BK006936.2| 513813 - INS 
 tpg|BK006947.3| 617995 + tpg|BK006947.3| 617641 - INS 
 tpg|BK006936.2| 645551 + tpg|BK006936.2| 645143 - INS 
 tpg|BK006947.3| 130339 + tpg|BK006947.3| 129784 - INS 
 tpg|BK006936.2| 789549 + tpg|BK006936.2| 788921 - INS 
 tpg|BK006947.3| 284485 + tpg|BK006947.3| 283880 - INS 
 tpg|BK006947.3| 628340 + tpg|BK006947.3| 628539 - INS 
 tpg|BK006936.2| 168657 + tpg|BK006936.2| 168028 - INS 
 tpg|BK006947.3| 537519 + tpg|BK006947.3| 537760 - INS 
 tpg|BK006947.3| 489609 + tpg|BK006947.3| 488861 - INS 
 tpg|BK006945.2| 727323 + tpg|BK006945.2| 726923 - INS 
 tpg|BK006947.3| 309333 + tpg|BK006947.3| 309064 - INS 
 tpg|BK006947.3| 509778 + tpg|BK006947.3| 510321 - INS 
 tpg|BK006945.2| 258790 + tpg|BK006945.2| 258492 - INS 
 tpg|BK006947.3| 185370 + tpg|BK006947.3| 185303 - INS 
 tpg|BK006945.2| 691279 + tpg|BK006945.2| 690600 - INS 
 tpg|BK006947.3| 220752 + tpg|BK006947.3| 220964 - INS 
 tpg|BK006947.3| 570181 + tpg|BK006947.3| 569870 - INS 
 tpg|BK006945.2| 680682 + tpg|BK006945.2| 681227 - INS 
 tpg|BK006947.3| 696648 + tpg|BK006947.3| 696333 - INS 
 tpg|BK006945.2| 420634 + tpg|BK006945.2| 419902 - INS 
 tpg|BK006947.3| 68191 + tpg|BK006947.3| 67721 - INS 
 tpg|BK006945.2| 417690 + tpg|BK006945.2| 417079 - INS 
 tpg|BK006945.2| 167295 + tpg|BK006945.2| 167580 - INS 
 tpg|BK006936.2| 775765 + tpg|BK006936.2| 775656 - INS 
 tpg|BK006945.2| 659382 + tpg|BK006945.2| 659791 - INS 
 tpg|BK006947.3| 753723 + tpg|BK006947.3| 754215 - INS 
 tpg|BK006947.3| 396435 + tpg|BK006947.3| 396288 - INS 
 tpg|BK006947.3| 393362 + tpg|BK006947.3| 392730 - INS 
 tpg|BK006945.2| 1041012 + tpg|BK006945.2| 1040855 - INS 
 tpg|BK006947.3| 295637 + tpg|BK006947.3| 295271 - INS 
 tpg|BK006936.2| 134745 + tpg|BK006936.2| 135162 - INS 
 tpg|BK006947.3| 336780 + tpg|BK006947.3| 336306 - INS 
 tpg|BK006947.3| 721507 + tpg|BK006947.3| 721071 - INS 
 tpg|BK006945.2| 381611 + tpg|BK006945.2| 381318 - INS 
 tpg|BK006936.2| 612900 + tpg|BK006936.2| 612863 - INS 
 tpg|BK006936.2| 698717 + tpg|BK006936.2| 699164 - INS 
 tpg|BK006947.3| 664413 + tpg|BK006947.3| 664328 - INS 
 tpg|BK006947.3| 55122 + tpg|BK006947.3| 54373 - INS 
 tpg|BK006947.3| 110569 + tpg|BK006947.3| 110038 - INS 
 tpg|BK006936.2| 456371 + tpg|BK006936.2| 456029 - INS 
 tpg|BK006947.3| 405716 + tpg|BK006947.3| 405679 - INS 
 tpg|BK006945.2| 576686 + tpg|BK006945.2| 577216 - INS 
 tpg|BK006947.3| 654640 + tpg|BK006947.3| 654393 - INS 
 tpg|BK006936.2| 449038 + tpg|BK006936.2| 448639 - INS 
 tpg|BK006947.3| 200127 + tpg|BK006947.3| 199526 - INS 
 tpg|BK006947.3| 399852 + tpg|BK006947.3| 400418 - INS 
 tpg|BK006936.2| 104230 + tpg|BK006936.2| 103647 - INS 
 tpg|BK006945.2| 104719 + tpg|BK006945.2| 104844 - INS 
 tpg|BK006947.3| 114174 + tpg|BK006947.3| 114059 - INS 
 tpg|BK006947.3| 370556 + tpg|BK006947.3| 369967 - INS 
 tpg|BK006936.2| 441624 + tpg|BK006936.2| 442173 - INS 
 tpg|BK006945.2| 29244 + tpg|BK006945.2| 28528 - INS 
 tpg|BK006947.3| 260267 + tpg|BK006947.3| 259957 - INS 
 tpg|BK006936.2| 544166 + tpg|BK006936.2| 543770 - INS A
 tpg|BK006947.3| 588962 + tpg|BK006947.3| 588420 - INS 
 tpg|BK006936.2| 420283 + tpg|BK006936.2| 420905 - INS 
 tpg|BK006947.3| 589659 + tpg|BK006947.3| 589154 - INS 
 tpg|BK006947.3| 341526 + tpg|BK006947.3| 341210 - INS 
 tpg|BK006947.3| 598087 + tpg|BK006947.3| 597672 - INS 
 tpg|BK006936.2| 454125 + tpg|BK006936.2| 454551 - INS 
 tpg|BK006947.3| 349227 + tpg|BK006947.3| 348462 - INS 
 tpg|BK006936.2| 556498 + tpg|BK006936.2| 556143 - INS 
 tpg|BK006947.3| 360968 + tpg|BK006947.3| 361401 - INS 
 tpg|BK006936.2| 292273 + tpg|BK006936.2| 291642 - INS 
 tpg|BK006947.3| 360038 + tpg|BK006947.3| 359435 - INS 
 tpg|BK006936.2| 293330 + tpg|BK006936.2| 293024 - INS 
 tpg|BK006936.2| 269500 + tpg|BK006936.2| 269903 - INS 
 tpg|BK006945.2| 322311 + tpg|BK006945.2| 322189 - INS 
 tpg|BK006947.3| 83807 + tpg|BK006947.3| 83513 - INS 
 tpg|BK006945.2| 511148 + tpg|BK006945.2| 511803 - INS 
 tpg|BK006936.2| 624553 + tpg|BK006936.2| 624348 - INS 
 tpg|BK006947.3| 774342 + tpg|BK006947.3| 774121 - INS 
 tpg|BK006945.2| 819797 + tpg|BK006945.2| 819627 - INS 
 tpg|BK006947.3| 685316 + tpg|BK006947.3| 685821 - INS 
 tpg|BK006936.2| 196240 + tpg|BK006936.2| 195705 - INS 
 tpg|BK006947.3| 597387 + tpg|BK006947.3| 596966 - INS 
 tpg|BK006947.3| 596459 + tpg|BK006947.3| 596589 - INS 
 tpg|BK006947.3| 694071 + tpg|BK006947.3| 693665 - INS 
 tpg|BK006947.3| 591599 + tpg|BK006947.3| 591490 - INS 
 tpg|BK006947.3| 496076 + tpg|BK006947.3| 495632 - INS 
 tpg|BK006947.3| 655536 + tpg|BK006947.3| 656113 - INS 
 tpg|BK006947.3| 190127 + tpg|BK006947.3| 189604 - INS 
 tpg|BK006936.2| 515593 + tpg|BK006936.2| 514914 - INS 
 tpg|BK006936.2| 724163 + tpg|BK006936.2| 723819 - INS 
 tpg|BK006947.3| 460271 + tpg|BK006947.3| 459795 - INS 
 tpg|BK006936.2| 722811 + tpg|BK006936.2| 722582 - INS 
 tpg|BK006947.3| 135547 + tpg|BK006947.3| 135355 - INS 
 tpg|BK006947.3| 235081 + tpg|BK006947.3| 234579 - INS 
 tpg|BK006936.2| 416938 + tpg|BK006936.2| 416887 - INS 
 tpg|BK006936.2| 12614 + tpg|BK006936.2| 12136 - INS 
 tpg|BK006947.3| 18347 + tpg|BK006947.3| 18656 - INS 
 tpg|BK006936.2| 70975 + tpg|BK006936.2| 71473 - INS 
 tpg|BK006947.3| 312709 + tpg|BK006947.3| 312192 - INS 
 tpg|BK006945.2| 489867 + tpg|BK006945.2| 489431 - INS 
 tpg|BK006936.2| 63977 + tpg|BK006936.2| 63631 - INS 
 tpg|BK006947.3| 652087 + tpg|BK006947.3| 651910 - INS 
 tpg|BK006945.2| 983553 + tpg|BK006945.2| 982857 - INS 
 tpg|BK006936.2| 52302 + tpg|BK006936.2| 51660 - INS 
 tpg|BK006947.3| 666974 + tpg|BK006947.3| 667135 - INS 
 tpg|BK006947.3| 325494 + tpg|BK006947.3| 326026 - INS TGG
 tpg|BK006936.2| 51129 + tpg|BK006936.2| 50870 - INS 
 tpg|BK006947.3| 104039 + tpg|BK006947.3| 104069 - INS 
 tpg|BK006945.2| 252689 + tpg|BK006945.2| 253290 - INS 
 tpg|BK006947.3| 218805 + tpg|BK006947.3| 218710 - INS 
 tpg|BK006936.2| 714181 + tpg|BK006936.2| 713434 - INS 
 tpg|BK006947.3| 254342 + tpg|BK006947.3| 254504 - INS 
 tpg|BK006936.2| 798435 + tpg|BK006936.2| 798608 - INS 
 tpg|BK006945.2| 272358 + tpg|BK006945.2| 272668 - INS 
 tpg|BK006947.3| 246522 + tpg|BK006947.3| 246457 - INS 
 tpg|BK006945.2| 1060265 + tpg|BK006945.2| 1059746 - INS 
 tpg|BK006947.3| 64500 + tpg|BK006947.3| 64195 - INS 
 tpg|BK006947.3| 233208 + tpg|BK006947.3| 233723 - INS 
 tpg|BK006936.2| 295530 + tpg|BK006936.2| 296086 - INS 
 tpg|BK006945.2| 622660 + tpg|BK006945.2| 622344 - INS 
 tpg|BK006947.3| 698594 + tpg|BK006947.3| 698537 - INS 
 tpg|BK006947.3| 235530 + tpg|BK006947.3| 235279 - INS 
 tpg|BK006947.3| 335004 + tpg|BK006947.3| 335324 - INS 
 tpg|BK006936.2| 357473 + tpg|BK006936.2| 356904 - INS 
 tpg|BK006936.2| 347399 + tpg|BK006936.2| 347816 - INS 
 tpg|BK006947.3| 557915 + tpg|BK006947.3| 557408 - INS 
 tpg|BK006947.3| 213551 + tpg|BK006947.3| 214133 - INS 
 tpg|BK006936.2| 123744 + tpg|BK006936.2| 123231 - INS 
 tpg|BK006947.3| 340237 + tpg|BK006947.3| 339837 - INS 
 tpg|BK006936.2| 490601 + tpg|BK006936.2| 490712 - INS 
 tpg|BK006947.3| 266591 + tpg|BK006947.3| 267182 - INS 
 tpg|BK006936.2| 581594 + tpg|BK006936.2| 581947 - INS 
 tpg|BK006947.3| 208298 + tpg|BK006947.3| 208114 - INS 
 tpg|BK006947.3| 500998 + tpg|BK006947.3| 501385 - INS 
 tpg|BK006936.2| 773189 + tpg|BK006936.2| 772740 - INS 
 tpg|BK006936.2| 258012 + tpg|BK006936.2| 257857 - INS 
 tpg|BK006945.2| 657310 + tpg|BK006945.2| 657050 - INS 
 tpg|BK006947.3| 552542 + tpg|BK006947.3| 551971 - INS 
 tpg|BK006947.3| 452393 + tpg|BK006947.3| 451729 - INS 
 tpg|BK006936.2| 441101 + tpg|BK006936.2| 441040 - INS 
 tpg|BK006936.2| 609214 + tpg|BK006936.2| 609385 - INS 
 tpg|BK006947.3| 32927 + tpg|BK006947.3| 32826 - INS 
 tpg|BK006936.2| 217787 + tpg|BK006936.2| 217096 - INS 
 tpg|BK006947.3| 587427 + tpg|BK006947.3| 587189 - INS 
 tpg|BK006936.2| 501398 + tpg|BK006936.2| 500948 - INS 
 tpg|BK006947.3| 368572 + tpg|BK006947.3| 367814 - INS 
 tpg|BK006947.3| 604098 + tpg|BK006947.3| 603810 - INS 
 tpg|BK006947.3| 61477 + tpg|BK006947.3| 60937 - INS 
 tpg|BK006936.2| 157577 + tpg|BK006936.2| 156820 - INS 
 tpg|BK006947.3| 28626 + tpg|BK006947.3| 27892 - INS 
 tpg|BK006947.3| 310730 + tpg|BK006947.3| 310575 - INS 
 tpg|BK006936.2| 142430 + tpg|BK006936.2| 143106 - INS 
 tpg|BK006936.2| 483213 + tpg|BK006936.2| 482798 - INS 
 tpg|BK006947.3| 536568 + tpg|BK006947.3| 536353 - INS 
 tpg|BK006947.3| 136293 + tpg|BK006947.3| 135972 - INS 
 tpg|BK006947.3| 186367 + tpg|BK006947.3| 186751 - INS 
 tpg|BK006945.2| 786764 + tpg|BK006945.2| 787455 - INS 
 tpg|BK006936.2| 662244 + tpg|BK006936.2| 661878 - INS 
 tpg|BK006947.3| 371456 + tpg|BK006947.3| 371697 - INS 
 tpg|BK006936.2| 125878 + tpg|BK006936.2| 125570 - INS 
 tpg|BK006947.3| 739157 + tpg|BK006947.3| 738406 - INS 
 tpg|BK006947.3| 412036 + tpg|BK006947.3| 411808 - INS 
 tpg|BK006945.2| 607037 + tpg|BK006945.2| 606887 - INS 
 tpg|BK006947.3| 204829 + tpg|BK006947.3| 204463 - INS 
 tpg|BK006947.3| 553531 + tpg|BK006947.3| 553576 - INS 
 tpg|BK006945.2| 229798 + tpg|BK006945.2| 229031 - INS 
 tpg|BK006947.3| 571345 + tpg|BK006947.3| 571980 - INS 
 tpg|BK006936.2| 105005 + tpg|BK006936.2| 104642 - INS 
 tpg|BK006945.2| 589472 + tpg|BK006945.2| 589331 - INS 
 tpg|BK006947.3| 572835 + tpg|BK006947.3| 572594 - INS 
 tpg|BK006947.3| 66931 + tpg|BK006947.3| 67288 - INS 
 tpg|BK006936.2| 122397 + tpg|BK006936.2| 121769 - INS 
 tpg|BK006947.3| 601304 + tpg|BK006947.3| 600857 - INS 
 tpg|BK006945.2| 926228 + tpg|BK006945.2| 925894 - INS 
 tpg|BK006947.3| 345426 + tpg|BK006947.3| 345457 - INS 
 tpg|BK006936.2| 523387 + tpg|BK006936.2| 523305 - INS 
 tpg|BK006947.3| 48656 + tpg|BK006947.3| 48640 - INS 
 tpg|BK006945.2| 397104 + tpg|BK006945.2| 396825 - INS 
 tpg|BK006947.3| 577538 + tpg|BK006947.3| 577882 - INS 
 tpg|BK006947.3| 303030 + tpg|BK006947.3| 303373 - INS 
 tpg|BK006936.2| 172521 + tpg|BK006936.2| 172876 - INS 
 tpg|BK006947.3| 485497 + tpg|BK006947.3| 484782 - INS 
 tpg|BK006936.2| 496447 + tpg|BK006936.2| 495846 - INS 
 tpg|BK006947.3| 211007 + tpg|BK006947.3| 210926 - INS 
 tpg|BK006936.2| 779969 + tpg|BK006936.2| 779757 - INS 
 tpg|BK006945.2| 120902 + tpg|BK006945.2| 120407 - INS 
 tpg|BK006947.3| 287487 + tpg|BK006947.3| 287121 - INS 
 tpg|BK006936.2| 679254 + tpg|BK006936.2| 678643 - INS 
 tpg|BK006947.3| 621028 + tpg|BK006947.3| 620789 - INS 
 tpg|BK006945.2| 89810 + tpg|BK006945.2| 89036 - INS 
 tpg|BK006947.3| 236614 + tpg|BK006947.3| 237064 - INS 
 tpg|BK006947.3| 602606 + tpg|BK006947.3| 601946 - INS 
 tpg|BK006947.3| 250828 + tpg|BK006947.3| 250728 - INS 
 tpg|BK006947.3| 682824 + tpg|BK006947.3| 682644 - INS 
 tpg|BK006936.2| 380910 + tpg|BK006936.2| 380683 - INS 
 tpg|BK006947.3| 677078 + tpg|BK006947.3| 677410 - INS 
 tpg|BK006947.3| 625382 + tpg|BK006947.3| 625033 - INS 
 tpg|BK006947.3| 257654 + tpg|BK006947.3| 257018 - INS 
 tpg|BK006936.2| 589382 + tpg|BK006936.2| 589674 - INS 
 tpg|BK006947.3| 280947 + tpg|BK006947.3| 280571 - INS 
 tpg|BK006947.3| 274737 + tpg|BK006947.3| 274246 - INS 
 tpg|BK006936.2| 458913 + tpg|BK006936.2| 458160 - INS 
 tpg|BK006947.3| 27080 + tpg|BK006947.3| 26759 - INS 
 tpg|BK006945.2| 829296 + tpg|BK006945.2| 828843 - INS 
 tpg|BK006947.3| 472559 + tpg|BK006947.3| 472891 - INS 
 tpg|BK006936.2| 592902 + tpg|BK006936.2| 592245 - INS 
 tpg|BK006947.3| 673603 + tpg|BK006947.3| 673399 - INS 
 tpg|BK006936.2| 321042 + tpg|BK006936.2| 320603 - INS 
 tpg|BK006947.3| 112130 + tpg|BK006947.3| 111687 - INS 
 tpg|BK006945.2| 200100 + tpg|BK006945.2| 199955 - INS 
 tpg|BK006947.3| 376599 + tpg|BK006947.3| 376906 - INS 
 tpg|BK006947.3| 474529 + tpg|BK006947.3| 474458 - INS 
 tpg|BK006945.2| 877913 + tpg|BK006945.2| 877679 - INS 
 tpg|BK006947.3| 366425 + tpg|BK006947.3| 365968 - INS 
 tpg|BK006947.3| 717582 + tpg|BK006947.3| 717249 - INS 
 tpg|BK006945.2| 939383 + tpg|BK006945.2| 940083 - INS 
 tpg|BK006947.3| 353615 + tpg|BK006947.3| 353497 - INS 
 tpg|BK006936.2| 805046 + tpg|BK006936.2| 804422 - INS 
 tpg|BK006947.3| 530473 + tpg|BK006947.3| 530431 - INS 
 tpg|BK006945.2| 601158 + tpg|BK006945.2| 601591 - INS 
 tpg|BK006936.2| 703469 + tpg|BK006936.2| 703385 - INS 
 tpg|BK006947.3| 523794 + tpg|BK006947.3| 523539 - INS 
 tpg|BK006945.2| 521737 + tpg|BK006945.2| 521357 - INS 
 tpg|BK006936.2| 23960 + tpg|BK006936.2| 24351 - INS 
 tpg|BK006947.3| 388268 + tpg|BK006947.3| 387901 - INS 
 tpg|BK006947.3| 670290 + tpg|BK006947.3| 670221 - INS 
 tpg|BK006936.2| 493976 + tpg|BK006936.2| 493477 - INS 
 tpg|BK006947.3| 681974 + tpg|BK006947.3| 681903 - INS 
 tpg|BK006947.3| 277537 + tpg|BK006947.3| 278295 - INS 
 tpg|BK006947.3| 410926 + tpg|BK006947.3| 410837 - INS 
 tpg|BK006936.2| 74817 + tpg|BK006936.2| 74054 - INS 
 tpg|BK006947.3| 151482 + tpg|BK006947.3| 151301 - INS 
 tpg|BK006945.2| 390210 + tpg|BK006945.2| 390527 - INS 
 tpg|BK006947.3| 150745 + tpg|BK006947.3| 150582 - INS 
 tpg|BK006936.2| 68073 + tpg|BK006936.2| 68163 - INS 
 tpg|BK006936.2| 182250 + tpg|BK006936.2| 182236 - INS 
 tpg|BK006947.3| 20658 + tpg|BK006947.3| 20484 - INS 
 tpg|BK006945.2| 524780 + tpg|BK006945.2| 524417 - INS 
 tpg|BK006936.2| 438799 + tpg|BK006936.2| 438613 - INS 
 tpg|BK006947.3| 313223 + tpg|BK006947.3| 313433 - INS 
 tpg|BK006947.3| 248720 + tpg|BK006947.3| 248455 - INS 
 tpg|BK006947.3| 154120 + tpg|BK006947.3| 153981 - INS 
 tpg|BK006945.2| 239376 + tpg|BK006945.2| 239837 - INS 
 tpg|BK006936.2| 304891 + tpg|BK006936.2| 304400 - INS 
 tpg|BK006947.3| 544530 + tpg|BK006947.3| 544114 - INS 
 tpg|BK006945.2| 262282 + tpg|BK006945.2| 262198 - INS 
 tpg|BK006947.3| 659234 + tpg|BK006947.3| 659115 - INS 
 tpg|BK006947.3| 539634 + tpg|BK006947.3| 539998 - INS 
 tpg|BK006947.3| 773419 + tpg|BK006947.3| 773057 - INS 
 tpg|BK006947.3| 176391 + tpg|BK006947.3| 176391 - INS 
 tpg|BK006945.2| 621040 + tpg|BK006945.2| 620994 - INS 
 tpg|BK006947.3| 611881 + tpg|BK006947.3| 611832 - INS 
 tpg|BK006947.3| 340910 + tpg|BK006947.3| 340614 - INS 
 tpg|BK006945.2| 520025 + tpg|BK006945.2| 519589 - INS 
 tpg|BK006947.3| 559168 + tpg|BK006947.3| 558484 - INS 
 tpg|BK006947.3| 609520 + tpg|BK006947.3| 609432 - INS 
 tpg|BK006947.3| 236208 + tpg|BK006947.3| 236051 - INS 
 tpg|BK006945.2| 230429 + tpg|BK006945.2| 229794 - INS 
 tpg|BK006947.3| 568972 + tpg|BK006947.3| 568802 - INS 
 tpg|BK006947.3| 222583 + tpg|BK006947.3| 222621 - INS 
 tpg|BK006945.2| 232966 + tpg|BK006945.2| 232757 - INS 
 tpg|BK006947.3| 245524 + tpg|BK006947.3| 244974 - INS 
 tpg|BK006945.2| 801971 + tpg|BK006945.2| 802489 - INS 
 tpg|BK006947.3| 759922 + tpg|BK006947.3| 759863 - INS 
 tpg|BK006945.2| 240039 + tpg|BK006945.2| 240381 - INS 
 tpg|BK006936.2| 607399 + tpg|BK006936.2| 607878 - INS 
 tpg|BK006947.3| 58532 + tpg|BK006947.3| 58355 - INS 
 tpg|BK006947.3| 101592 + tpg|BK006947.3| 101422 - INS 
 tpg|BK006945.2| 918568 + tpg|BK006945.2| 917924 - INS 
 tpg|BK006947.3| 558400 + tpg|BK006947.3| 557847 - INS 
 tpg|BK006947.3| 255355 + tpg|BK006947.3| 255877 - INS 
 tpg|BK006947.3| 414621 + tpg|BK006947.3| 414548 - INS 
 tpg|BK006947.3| 110968 + tpg|BK006947.3| 111066 - INS 
 tpg|BK006947.3| 467985 + tpg|BK006947.3| 468510 - INS 
 tpg|BK006947.3| 382258 + tpg|BK006947.3| 381669 - INS 
 tpg|BK006947.3| 360345 + tpg|BK006947.3| 360467 - INS 
 tpg|BK006947.3| 764030 + tpg|BK006947.3| 764439 - INS 
 tpg|BK006947.3| 436864 + tpg|BK006947.3| 437000 - INS 
 tpg|BK006945.2| 638933 + tpg|BK006945.2| 638384 - INS 
 tpg|BK006947.3| 269472 + tpg|BK006947.3| 268987 - INS 
 tpg|BK006947.3| 318511 + tpg|BK006947.3| 318418 - INS 
 tpg|BK006947.3| 154448 + tpg|BK006947.3| 155189 - INS 
 tpg|BK006947.3| 443146 + tpg|BK006947.3| 443235 - INS 
 tpg|BK006945.2| 1013344 + tpg|BK006945.2| 1014093 - INS 
 tpg|BK006947.3| 136958 + tpg|BK006947.3| 136679 - INS 
 tpg|BK006947.3| 647384 + tpg|BK006947.3| 647358 - INS 
 tpg|BK006947.3| 258196 + tpg|BK006947.3| 258737 - INS 
 tpg|BK006947.3| 545031 + tpg|BK006947.3| 544730 - INS 
 tpg|BK006945.2| 118808 + tpg|BK006945.2| 118242 - INS 
 tpg|BK006947.3| 438663 + tpg|BK006947.3| 437910 - INS 
 tpg|BK006947.3| 390570 + tpg|BK006947.3| 390416 - INS 
 tpg|BK006947.3| 496443 + tpg|BK006947.3| 496495 - INS 
 tpg|BK006945.2| 993601 + tpg|BK006945.2| 992900 - INS 
 tpg|BK006947.3| 369085 + tpg|BK006947.3| 368624 - INS 
 tpg|BK006947.3| 165913 + tpg|BK006947.3| 165593 - INS 
 tpg|BK006945.2| 874748 + tpg|BK006945.2| 874717 - INS 
 tpg|BK006947.3| 539178 + tpg|BK006947.3| 538789 - INS 
 tpg|BK006945.2| 935429 + tpg|BK006945.2| 934817 - INS 
 tpg|BK006947.3| 280241 + tpg|BK006947.3| 280082 - INS 
 tpg|BK006947.3| 775199 + tpg|BK006947.3| 774874 - INS 
 tpg|BK006947.3| 579824 + tpg|BK006947.3| 580484 - INS 
 tpg|BK006947.3| 606759 + tpg|BK006947.3| 606598 - INS 
 tpg|BK006945.2| 997907 + tpg|BK006945.2| 997892 - INS 
 tpg|BK006945.2| 996998 + tpg|BK006945.2| 996745 - INS 
 tpg|BK006945.2| 541600 + tpg|BK006945.2| 540857 - INS 
 tpg|BK006945.2| 605509 + tpg|BK006945.2| 605979 - INS 
 tpg|BK006945.2| 704163 + tpg|BK006945.2| 703647 - INS 
 tpg|BK006945.2| 441940 + tpg|BK006945.2| 442331 - INS 
 tpg|BK006945.2| 812730 + tpg|BK006945.2| 812026 - INS 
 tpg|BK006945.2| 301846 + tpg|BK006945.2| 301997 - INS 
 tpg|BK006945.2| 429409 + tpg|BK006945.2| 429866 - INS 
 tpg|BK006945.2| 677153 + tpg|BK006945.2| 676490 - INS 
 tpg|BK006945.2| 773447 + tpg|BK006945.2| 773177 - INS 
 tpg|BK006945.2| 450347 + tpg|BK006945.2| 449984 - INS 
 tpg|BK006945.2| 760202 + tpg|BK006945.2| 760333 - INS 
 tpg|BK006945.2| 34191 + tpg|BK006945.2| 34693 - INS 
 tpg|BK006945.2| 221896 + tpg|BK006945.2| 222178 - INS 
 tpg|BK006945.2| 824642 + tpg|BK006945.2| 824579 - INS 
 tpg|BK006945.2| 371463 + tpg|BK006945.2| 370985 - INS 
 tpg|BK006945.2| 376600 + tpg|BK006945.2| 376663 - INS 
 tpg|BK006945.2| 1038861 + tpg|BK006945.2| 1039454 - INS 
 tpg|BK006945.2| 425519 + tpg|BK006945.2| 425239 - INS 
 tpg|BK006945.2| 351412 + tpg|BK006945.2| 350697 - INS 
 tpg|BK006945.2| 785626 + tpg|BK006945.2| 785682 - INS 
 tpg|BK006945.2| 328908 + tpg|BK006945.2| 328476 - INS 
 tpg|BK006945.2| 827356 + tpg|BK006945.2| 827060 - INS 
 tpg|BK006945.2| 364794 + tpg|BK006945.2| 364366 - INS 
 tpg|BK006945.2| 413112 + tpg|BK006945.2| 413147 - INS 
 tpg|BK006945.2| 983886 + tpg|BK006945.2| 983542 - INS 
 tpg|BK006945.2| 116725 + tpg|BK006945.2| 116949 - INS 
 tpg|BK006945.2| 255167 + tpg|BK006945.2| 254929 - INS 
 tpg|BK006945.2| 562184 + tpg|BK006945.2| 562019 - INS 
 tpg|BK006945.2| 241402 + tpg|BK006945.2| 241480 - INS 
 tpg|BK006936.2| 1965 + tpg|BK006936.2| 1729 - INS CTAG
 tpg|BK006936.2| 466741 + tpg|BK006936.2| 466023 - INS 
 tpg|BK006936.2| 739369 + tpg|BK006936.2| 739777 - INS 
 tpg|BK006936.2| 410077 + tpg|BK006936.2| 410362 - INS 
 tpg|BK006936.2| 808755 + tpg|BK006936.2| 808070 - INS 
 tpg|BK006936.2| 475240 + tpg|BK006936.2| 474719 - INS 
 tpg|BK006936.2| 322232 + tpg|BK006936.2| 322721 - INS 
 tpg|BK006936.2| 16714 + tpg|BK006936.2| 16477 - INS 
 tpg|BK006936.2| 218305 + tpg|BK006936.2| 217967 - INS 
 tpg|BK006936.2| 268785 + tpg|BK006936.2| 269213 - INS 
 tpg|BK006936.2| 683133 + tpg|BK006936.2| 682719 - INS 
 tpg|BK006936.2| 488846 + tpg|BK006936.2| 489004 - INS 
 tpg|BK006936.2| 582063 + tpg|BK006936.2| 582480 - INS 
 tpg|BK006936.2| 319419 + tpg|BK006936.2| 319821 - INS 
 tpg|BK006936.2| 800367 + tpg|BK006936.2| 801060 - INS 
 tpg|BK006936.2| 251938 + tpg|BK006936.2| 251197 - INS 
 tpg|BK006936.2| 245172 + tpg|BK006936.2| 244660 - INS 
 tpg|BK006936.2| 330799 + tpg|BK006936.2| 330182 - INS 
 tpg|BK006936.2| 307898 + tpg|BK006936.2| 307688 - INS 
 tpg|BK006936.2| 665412 + tpg|BK006936.2| 665301 - INS 
 tpg|BK006936.2| 632589 + tpg|BK006936.2| 632271 - INS 
 tpg|BK006936.2| 633968 + tpg|BK006936.2| 634011 - INS 
 tpg|BK006936.2| 192320 + tpg|BK006936.2| 192132 - INS 
 tpg|BK006936.2| 524714 + tpg|BK006936.2| 524429 - INS 
 tpg|BK006936.2| 174367 + tpg|BK006936.2| 173855 - INS 
 tpg|BK006936.2| 154760 + tpg|BK006936.2| 154911 - INS 
 tpg|BK006936.2| 781065 + tpg|BK006936.2| 781356 - INS 
 tpg|BK006936.2| 378517 + tpg|BK006936.2| 377888 - INS 
 tpg|BK006936.2| 187333 + tpg|BK006936.2| 187675 - INS 
 tpg|BK006936.2| 189945 + tpg|BK006936.2| 189701 - INS 
 tpg|BK006936.2| 668786 + tpg|BK006936.2| 668902 - INS 
 tpg|BK006936.2| 327048 + tpg|BK006936.2| 326728 - INS 
 tpg|BK006936.2| 151938 + tpg|BK006936.2| 151644 - INS 
 tpg|BK006936.2| 435247 + tpg|BK006936.2| 435267 - INS 
 tpg|BK006936.2| 603785 + tpg|BK006936.2| 603897 - INS 
 tpg|BK006936.2| 741032 + tpg|BK006936.2| 741387 - INS 
 tpg|BK006936.2| 362293 + tpg|BK006936.2| 362981 - INS 
 tpg|BK006936.2| 506387 + tpg|BK006936.2| 506299 - INS 
 tpg|BK006936.2| 154043 + tpg|BK006936.2| 153321 - INS 
 tpg|BK006936.2| 361466 + tpg|BK006936.2| 360794 - INS 
 tpg|BK006936.2| 215524 + tpg|BK006936.2| 215352 - INS 
 tpg|BK006936.2| 577473 + tpg|BK006936.2| 577310 - INS 
 tpg|BK006936.2| 287264 + tpg|BK006936.2| 287738 - INS 
 tpg|BK006936.2| 507889 + tpg|BK006936.2| 507931 - INS 
 tpg|BK006936.2| 720293 + tpg|BK006936.2| 720129 - INS 
 tpg|BK006936.2| 400399 + tpg|BK006936.2| 400048 - INS 
 tpg|BK006936.2| 42816 + tpg|BK006936.2| 43452 - INS 
 tpg|BK006936.2| 101248 + tpg|BK006936.2| 100729 - INS 
 tpg|BK006936.2| 180430 + tpg|BK006936.2| 180906 - INS 
 tpg|BK006936.2| 92280 + tpg|BK006936.2| 91571 - INS 
 tpg|BK006945.2| 903086 + tpg|BK006945.2| 902676 - INS 
 tpg|BK006936.2| 411193 + tpg|BK006936.2| 411273 - INS 
 tpg|BK006945.2| 395618 + tpg|BK006945.2| 395169 - INS 
 tpg|BK006936.2| 58695 + tpg|BK006936.2| 58994 - INS 
 tpg|BK006945.2| 339885 + tpg|BK006945.2| 339744 - INS 
 tpg|BK006945.2| 723052 + tpg|BK006945.2| 722290 - INS 
 tpg|BK006945.2| 434594 + tpg|BK006945.2| 434448 - INS 
 tpg|BK006945.2| 106780 + tpg|BK006945.2| 107423 - INS 
 tpg|BK006945.2| 917531 + tpg|BK006945.2| 917132 - INS 
 tpg|BK006945.2| 251191 + tpg|BK006945.2| 250484 - INS 
 tpg|BK006936.2| 165927 + tpg|BK006936.2| 165911 - INS 
 tpg|BK006936.2| 11397 + tpg|BK006936.2| 11274 - INS 
 tpg|BK006945.2| 544222 + tpg|BK006945.2| 544451 - INS 
 tpg|BK006936.2| 486417 + tpg|BK006936.2| 486990 - INS 
 tpg|BK006945.2| 503749 + tpg|BK006945.2| 503874 - INS 
 tpg|BK006936.2| 387412 + tpg|BK006936.2| 386953 - INS 
 tpg|BK006936.2| 388473 + tpg|BK006936.2| 388272 - INS 
 tpg|BK006945.2| 347584 + tpg|BK006945.2| 347632 - INS 
 tpg|BK006945.2| 208060 + tpg|BK006945.2| 208158 - INS 
 tpg|BK006936.2| 389598 + tpg|BK006936.2| 389115 - INS 
 tpg|BK006936.2| 712774 + tpg|BK006936.2| 712498 - INS 
 tpg|BK006936.2| 101759 + tpg|BK006936.2| 101966 - INS 
 tpg|BK006936.2| 406156 + tpg|BK006936.2| 406500 - INS 
 tpg|BK006945.2| 332921 + tpg|BK006945.2| 333365 - INS 
 tpg|BK006936.2| 737648 + tpg|BK006936.2| 737506 - INS 
 tpg|BK006936.2| 716989 + tpg|BK006936.2| 717017 - INS 
 tpg|BK006945.2| 865984 + tpg|BK006945.2| 865960 - INS 
 tpg|BK006936.2| 554302 + tpg|BK006936.2| 554969 - INS 
 tpg|BK006936.2| 287975 + tpg|BK006936.2| 288161 - INS 
 tpg|BK006945.2| 329622 + tpg|BK006945.2| 330057 - INS 
 tpg|BK006936.2| 562392 + tpg|BK006936.2| 563023 - INS 
 tpg|BK006936.2| 248030 + tpg|BK006936.2| 248183 - INS 
 tpg|BK006945.2| 311944 + tpg|BK006945.2| 312181 - INS 
 tpg|BK006936.2| 616247 + tpg|BK006936.2| 616392 - INS 
 tpg|BK006945.2| 120045 + tpg|BK006945.2| 119922 - INS 
 tpg|BK006936.2| 337507 + tpg|BK006936.2| 337405 - INS 
 tpg|BK006945.2| 292557 + tpg|BK006945.2| 291972 - INS 
 tpg|BK006945.2| 18492 + tpg|BK006945.2| 18427 - INS 
 tpg|BK006936.2| 516462 + tpg|BK006936.2| 516303 - INS 
 tpg|BK006936.2| 725377 + tpg|BK006936.2| 724977 - INS 
 tpg|BK006945.2| 537160 + tpg|BK006945.2| 537492 - INS 
 tpg|BK006936.2| 36966 + tpg|BK006936.2| 37282 - INS 
 tpg|BK006945.2| 110554 + tpg|BK006945.2| 110365 - INS 
 tpg|BK006945.2| 844043 + tpg|BK006945.2| 843479 - INS ACAA
 tpg|BK006936.2| 357838 + tpg|BK006936.2| 357375 - INS 
 tpg|BK006945.2| 70569 + tpg|BK006945.2| 69954 - INS 
 tpg|BK006945.2| 587744 + tpg|BK006945.2| 587472 - INS 
 tpg|BK006936.2| 672008 + tpg|BK006936.2| 672745 - INS 
 tpg|BK006936.2| 680759 + tpg|BK006936.2| 681004 - INS 
 tpg|BK006945.2| 15391 + tpg|BK006945.2| 15055 - INS 
 tpg|BK006936.2| 697589 + tpg|BK006936.2| 698154 - INS 
 tpg|BK006945.2| 571439 + tpg|BK006945.2| 570749 - INS 
 tpg|BK006936.2| 190707 + tpg|BK006936.2| 190888 - INS 
 tpg|BK006936.2| 801515 + tpg|BK006936.2| 801474 - INS 
 tpg|BK006936.2| 740584 + tpg|BK006936.2| 740326 - INS 
 tpg|BK006945.2| 542086 + tpg|BK006945.2| 541419 - INS 
 tpg|BK006945.2| 815309 + tpg|BK006945.2| 815714 - INS 
 tpg|BK006945.2| 530164 + tpg|BK006945.2| 529983 - INS 
 tpg|BK006945.2| 611563 + tpg|BK006945.2| 611277 - INS 
 tpg|BK006936.2| 239695 + tpg|BK006936.2| 240197 - INS GCTCCACCATA
 tpg|BK006936.2| 351311 + tpg|BK006936.2| 350688 - INS 
 tpg|BK006945.2| 95554 + tpg|BK006945.2| 95479 - INS 
 tpg|BK006945.2| 620129 + tpg|BK006945.2| 620067 - INS 
 tpg|BK006936.2| 674631 + tpg|BK006936.2| 675073 - INS 
 tpg|BK006945.2| 857230 + tpg|BK006945.2| 856539 - INS 
 tpg|BK006945.2| 491640 + tpg|BK006945.2| 491514 - INS 
 tpg|BK006936.2| 249048 + tpg|BK006936.2| 249092 - INS 
 tpg|BK006936.2| 599945 + tpg|BK006936.2| 600631 - INS 
 tpg|BK006945.2| 1044591 + tpg|BK006945.2| 1044121 - INS 
 tpg|BK006945.2| 674452 + tpg|BK006945.2| 673804 - INS 
 tpg|BK006936.2| 159296 + tpg|BK006936.2| 159664 - INS 
 tpg|BK006945.2| 62093 + tpg|BK006945.2| 61795 - INS 
 tpg|BK006936.2| 277426 + tpg|BK006936.2| 277196 - INS 
 tpg|BK006936.2| 280602 + tpg|BK006936.2| 280228 - INS 
 tpg|BK006936.2| 335443 + tpg|BK006936.2| 335535 - INS 
 tpg|BK006945.2| 159746 + tpg|BK006945.2| 159692 - INS CTA
 tpg|BK006936.2| 655576 + tpg|BK006936.2| 655812 - INS 
 tpg|BK006936.2| 282635 + tpg|BK006936.2| 281883 - INS 
 tpg|BK006945.2| 38827 + tpg|BK006945.2| 38247 - INS 
 tpg|BK006936.2| 485944 + tpg|BK006936.2| 485288 - INS 
 tpg|BK006945.2| 658269 + tpg|BK006945.2| 657923 - INS 
 tpg|BK006936.2| 427481 + tpg|BK006936.2| 427813 - INS 
 tpg|BK006945.2| 436180 + tpg|BK006945.2| 435628 - INS 
 tpg|BK006936.2| 397289 + tpg|BK006936.2| 397295 - INS 
 tpg|BK006945.2| 646395 + tpg|BK006945.2| 646391 - INS 
 tpg|BK006945.2| 394965 + tpg|BK006945.2| 394603 - INS 
 tpg|BK006936.2| 730960 + tpg|BK006936.2| 731532 - INS 
 tpg|BK006936.2| 88369 + tpg|BK006936.2| 87901 - INS 
 tpg|BK006945.2| 989084 + tpg|BK006945.2| 988723 - INS 
 tpg|BK006945.2| 643899 + tpg|BK006945.2| 643280 - INS 
 tpg|BK006936.2| 748338 + tpg|BK006936.2| 748092 - INS 
 tpg|BK006936.2| 426686 + tpg|BK006936.2| 426425 - INS 
 tpg|BK006936.2| 276019 + tpg|BK006936.2| 275648 - INS 
 tpg|BK006936.2| 26015 + tpg|BK006936.2| 26129 - INS 
 tpg|BK006936.2| 48015 + tpg|BK006936.2| 48123 - INS 
 tpg|BK006936.2| 332006 + tpg|BK006936.2| 331496 - INS 
 tpg|BK006936.2| 208605 + tpg|BK006936.2| 207899 - INS 
 tpg|BK006936.2| 202016 + tpg|BK006936.2| 201280 - INS 
 tpg|BK006936.2| 689501 + tpg|BK006936.2| 689744 - INS 
 tpg|BK006945.2| 374655 + tpg|BK006945.2| 374826 - INS 
 tpg|BK006936.2| 353229 + tpg|BK006936.2| 352585 - INS 
 tpg|BK006945.2| 378096 + tpg|BK006945.2| 377547 - INS 
 tpg|BK006936.2| 354543 + tpg|BK006936.2| 354245 - INS 
 tpg|BK006945.2| 93272 + tpg|BK006945.2| 92874 - INS 
 tpg|BK006945.2| 689843 + tpg|BK006945.2| 689336 - INS 
 tpg|BK006936.2| 704824 + tpg|BK006936.2| 704149 - INS 
 tpg|BK006945.2| 700626 + tpg|BK006945.2| 699970 - INS 
 tpg|BK006936.2| 705358 + tpg|BK006936.2| 705239 - INS 
 tpg|BK006936.2| 231563 + tpg|BK006936.2| 232258 - INS 
 tpg|BK006936.2| 652766 + tpg|BK006936.2| 653011 - INS 
 tpg|BK006945.2| 698979 + tpg|BK006945.2| 698811 - INS 
 tpg|BK006945.2| 386960 + tpg|BK006945.2| 386589 - INS 
 tpg|BK006936.2| 520105 + tpg|BK006936.2| 519894 - INS 
 tpg|BK006936.2| 202499 + tpg|BK006936.2| 202999 - INS 
 tpg|BK006936.2| 170219 + tpg|BK006936.2| 169926 - INS 
 tpg|BK006936.2| 671456 + tpg|BK006936.2| 671080 - INS 
 tpg|BK006936.2| 429535 + tpg|BK006936.2| 429141 - INS 
 tpg|BK006936.2| 14665 + tpg|BK006936.2| 14881 - INS 
 tpg|BK006945.2| 380120 + tpg|BK006945.2| 379487 - INS 
 tpg|BK006936.2| 674133 + tpg|BK006936.2| 673869 - INS 
 tpg|BK006945.2| 702901 + tpg|BK006945.2| 702660 - INS 
 tpg|BK006936.2| 792165 + tpg|BK006936.2| 791410 - INS 
 tpg|BK006936.2| 407806 + tpg|BK006936.2| 407056 - INS 
 tpg|BK006936.2| 42080 + tpg|BK006936.2| 41670 - INS 
 tpg|BK006936.2| 610369 + tpg|BK006936.2| 610138 - INS 
 tpg|BK006945.2| 67504 + tpg|BK006945.2| 67534 - INS 
 tpg|BK006945.2| 542901 + tpg|BK006945.2| 543019 - INS 
 tpg|BK006936.2| 381887 + tpg|BK006936.2| 381505 - INS 
 tpg|BK006936.2| 752898 + tpg|BK006936.2| 752690 - INS 
 tpg|BK006945.2| 921189 + tpg|BK006945.2| 921190 - INS 
 tpg|BK006936.2| 376679 + tpg|BK006936.2| 376140 - INS 
 tpg|BK006945.2| 539534 + tpg|BK006945.2| 539678 - INS 
 tpg|BK006936.2| 487667 + tpg|BK006936.2| 487931 - INS 
 tpg|BK006945.2| 873979 + tpg|BK006945.2| 873786 - INS 
 tpg|BK006936.2| 400831 + tpg|BK006936.2| 401357 - INS 
 tpg|BK006945.2| 871533 + tpg|BK006945.2| 870831 - INS 
 tpg|BK006936.2| 491585 + tpg|BK006936.2| 491897 - INS 
 tpg|BK006936.2| 306326 + tpg|BK006936.2| 306087 - INS 
 tpg|BK006945.2| 318079 + tpg|BK006945.2| 318316 - INS 
 tpg|BK006945.2| 1055571 + tpg|BK006945.2| 1054809 - INS 
 tpg|BK006936.2| 588352 + tpg|BK006936.2| 587813 - INS 
 tpg|BK006936.2| 715572 + tpg|BK006936.2| 715214 - INS 
 tpg|BK006936.2| 799459 + tpg|BK006936.2| 799278 - INS 
 tpg|BK006936.2| 450242 + tpg|BK006936.2| 449703 - INS 
 tpg|BK006936.2| 132571 + tpg|BK006936.2| 132303 - INS 
 tpg|BK006936.2| 334354 + tpg|BK006936.2| 334637 - INS 
 tpg|BK006945.2| 243016 + tpg|BK006945.2| 242485 - INS 
 tpg|BK006936.2| 677252 + tpg|BK006936.2| 677765 - INS 
 tpg|BK006936.2| 158445 + tpg|BK006936.2| 158342 - INS 
 tpg|BK006945.2| 627527 + tpg|BK006945.2| 627035 - INS 
 tpg|BK006945.2| 600288 + tpg|BK006945.2| 599575 - INS 
 tpg|BK006936.2| 536787 + tpg|BK006936.2| 537015 - INS 
 tpg|BK006945.2| 277770 + tpg|BK006945.2| 277881 - INS 
 tpg|BK006936.2| 652208 + tpg|BK006936.2| 651620 - INS 
 tpg|BK006936.2| 546556 + tpg|BK006936.2| 547103 - INS 
 tpg|BK006945.2| 189834 + tpg|BK006945.2| 189268 - INS 
 tpg|BK006936.2| 658166 + tpg|BK006936.2| 657481 - INS 
 tpg|BK006936.2| 284487 + tpg|BK006936.2| 285183 - INS 
 tpg|BK006945.2| 953422 + tpg|BK006945.2| 953481 - INS 
 tpg|BK006936.2| 221374 + tpg|BK006936.2| 220862 - INS 
 tpg|BK006945.2| 446721 + tpg|BK006945.2| 447318 - INS 
 tpg|BK006936.2| 614061 + tpg|BK006936.2| 614417 - INS 
 tpg|BK006945.2| 610484 + tpg|BK006945.2| 609933 - INS 
 tpg|BK006936.2| 591436 + tpg|BK006936.2| 590869 - INS 
 tpg|BK006945.2| 431788 + tpg|BK006945.2| 431370 - INS 
 tpg|BK006936.2| 638264 + tpg|BK006936.2| 638774 - INS 
 tpg|BK006936.2| 643440 + tpg|BK006936.2| 642720 - INS 
 tpg|BK006936.2| 637372 + tpg|BK006936.2| 636796 - INS 
 tpg|BK006936.2| 636567 + tpg|BK006936.2| 636212 - INS 
 tpg|BK006936.2| 242436 + tpg|BK006936.2| 241984 - INS 
 tpg|BK006945.2| 706535 + tpg|BK006945.2| 706223 - INS 
 tpg|BK006945.2| 369529 + tpg|BK006945.2| 369325 - INS 
 tpg|BK006936.2| 759439 + tpg|BK006936.2| 758876 - INS 
 tpg|BK006945.2| 771102 + tpg|BK006945.2| 771509 - INS 
 tpg|BK006945.2| 774923 + tpg|BK006945.2| 774577 - INS 
 tpg|BK006936.2| 759886 + tpg|BK006936.2| 759584 - INS 
 tpg|BK006936.2| 484061 + tpg|BK006936.2| 483409 - INS 
 tpg|BK006945.2| 102206 + tpg|BK006945.2| 102077 - INS 
 tpg|BK006945.2| 567927 + tpg|BK006945.2| 568023 - INS 
 tpg|BK006945.2| 719396 + tpg|BK006945.2| 720088 - INS 
 tpg|BK006936.2| 498821 + tpg|BK006936.2| 498510 - INS 
 tpg|BK006936.2| 80741 + tpg|BK006936.2| 80510 - INS 
 tpg|BK006945.2| 830626 + tpg|BK006945.2| 830744 - INS 
 tpg|BK006936.2| 757908 + tpg|BK006936.2| 757252 - INS 
 tpg|BK006936.2| 428675 + tpg|BK006936.2| 428449 - INS 
 tpg|BK006945.2| 569452 + tpg|BK006945.2| 570161 - INS 
 tpg|BK006936.2| 548947 + tpg|BK006936.2| 549230 - INS 
 tpg|BK006936.2| 431572 + tpg|BK006936.2| 431232 - INS 
 tpg|BK006945.2| 975521 + tpg|BK006945.2| 974792 - INS 
 tpg|BK006936.2| 358798 + tpg|BK006936.2| 359411 - INS 
 tpg|BK006945.2| 275619 + tpg|BK006945.2| 275990 - INS 
 tpg|BK006936.2| 644112 + tpg|BK006936.2| 644389 - INS 
 tpg|BK006945.2| 973558 + tpg|BK006945.2| 973427 - INS 
 tpg|BK006936.2| 90300 + tpg|BK006936.2| 90683 - INS 
 tpg|BK006936.2| 97374 + tpg|BK006936.2| 97924 - INS 
 tpg|BK006945.2| 249904 + tpg|BK006945.2| 249866 - INS 
 tpg|BK006936.2| 250357 + tpg|BK006936.2| 250114 - INS 
 tpg|BK006936.2| 598728 + tpg|BK006936.2| 598718 - INS 
 tpg|BK006936.2| 349087 + tpg|BK006936.2| 348990 - INS 
 tpg|BK006936.2| 126384 + tpg|BK006936.2| 126186 - INS 
 tpg|BK006936.2| 694455 + tpg|BK006936.2| 693794 - INS 
 tpg|BK006936.2| 150717 + tpg|BK006936.2| 151041 - INS 
 tpg|BK006936.2| 670771 + tpg|BK006936.2| 670042 - INS 
 tpg|BK006936.2| 663118 + tpg|BK006936.2| 662696 - INS 
 tpg|BK006936.2| 183262 + tpg|BK006936.2| 183446 - INS 
 tpg|BK006936.2| 54895 + tpg|BK006936.2| 55408 - INS 
 tpg|BK006945.2| 245537 + tpg|BK006945.2| 245713 - INS 
 tpg|BK006936.2| 186566 + tpg|BK006936.2| 186430 - INS 
 tpg|BK006936.2| 553231 + tpg|BK006936.2| 552941 - INS 
 tpg|BK006936.2| 201117 + tpg|BK006936.2| 200701 - INS 
 tpg|BK006945.2| 20456 + tpg|BK006945.2| 20309 - INS 
 tpg|BK006936.2| 737120 + tpg|BK006936.2| 736652 - INS 
 tpg|BK006936.2| 542496 + tpg|BK006936.2| 542362 - INS 
 tpg|BK006945.2| 523968 + tpg|BK006945.2| 523289 - INS 
 tpg|BK006936.2| 20887 + tpg|BK006936.2| 20149 - INS 
 tpg|BK006936.2| 171312 + tpg|BK006936.2| 171466 - INS 
 tpg|BK006945.2| 74928 + tpg|BK006945.2| 74568 - INS 
 tpg|BK006936.2| 242915 + tpg|BK006936.2| 243479 - INS 
 tpg|BK006936.2| 227618 + tpg|BK006936.2| 227924 - INS 
 tpg|BK006936.2| 178794 + tpg|BK006936.2| 178625 - INS 
 tpg|BK006945.2| 234020 + tpg|BK006945.2| 234604 - INS 
 tpg|BK006936.2| 109698 + tpg|BK006936.2| 109263 - INS 
 tpg|BK006936.2| 371258 + tpg|BK006936.2| 371430 - INS 
 tpg|BK006945.2| 25457 + tpg|BK006945.2| 24820 - INS 
 tpg|BK006936.2| 374739 + tpg|BK006936.2| 374540 - INS 
 tpg|BK006936.2| 219400 + tpg|BK006936.2| 218772 - INS 
 tpg|BK006936.2| 199664 + tpg|BK006936.2| 199792 - INS 
 tpg|BK006945.2| 130126 + tpg|BK006945.2| 130452 - INS 
 tpg|BK006936.2| 213732 + tpg|BK006936.2| 213248 - INS 
 tpg|BK006936.2| 377023 + tpg|BK006936.2| 376715 - INS 
 tpg|BK006936.2| 539619 + tpg|BK006936.2| 539204 - INS 
 tpg|BK006936.2| 382435 + tpg|BK006936.2| 381981 - INS 
 tpg|BK006936.2| 796070 + tpg|BK006936.2| 796267 - INS 
 tpg|BK006936.2| 148254 + tpg|BK006936.2| 147568 - INS 
 tpg|BK006936.2| 628024 + tpg|BK006936.2| 627698 - INS 
 tpg|BK006936.2| 484650 + tpg|BK006936.2| 484747 - INS 
 tpg|BK006945.2| 1049760 + tpg|BK006945.2| 1049721 - INS 
 tpg|BK006945.2| 314866 + tpg|BK006945.2| 314223 - INS 
 tpg|BK006936.2| 633054 + tpg|BK006936.2| 632735 - INS 
 tpg|BK006945.2| 88105 + tpg|BK006945.2| 87427 - INS 
 tpg|BK006936.2| 305691 + tpg|BK006936.2| 305411 - INS 
 tpg|BK006945.2| 144916 + tpg|BK006945.2| 144834 - INS 
 tpg|BK006936.2| 752381 + tpg|BK006936.2| 751838 - INS 
 tpg|BK006936.2| 138141 + tpg|BK006936.2| 137786 - INS 
 tpg|BK006945.2| 640974 + tpg|BK006945.2| 640997 - INS 
 tpg|BK006936.2| 197625 + tpg|BK006936.2| 197608 - INS 
 tpg|BK006936.2| 238740 + tpg|BK006936.2| 238313 - INS 
 tpg|BK006945.2| 336960 + tpg|BK006945.2| 336849 - INS 
 tpg|BK006945.2| 742672 + tpg|BK006945.2| 742474 - INS 
 tpg|BK006936.2| 339304 + tpg|BK006936.2| 338537 - INS 
 tpg|BK006936.2| 477349 + tpg|BK006936.2| 477104 - INS 
 tpg|BK006945.2| 214984 + tpg|BK006945.2| 214587 - INS 
 tpg|BK006936.2| 117804 + tpg|BK006936.2| 118255 - INS 
 tpg|BK006945.2| 878724 + tpg|BK006945.2| 879102 - INS 
 tpg|BK006936.2| 70351 + tpg|BK006936.2| 69962 - INS 
 tpg|BK006936.2| 283358 + tpg|BK006936.2| 282802 - INS 
 tpg|BK006936.2| 666352 + tpg|BK006936.2| 666893 - INS 
 tpg|BK006936.2| 323463 + tpg|BK006936.2| 323144 - INS 
 tpg|BK006936.2| 163455 + tpg|BK006936.2| 163817 - INS 
 tpg|BK006945.2| 576056 + tpg|BK006945.2| 576717 - INS 
 tpg|BK006936.2| 351785 + tpg|BK006936.2| 351326 - INS 
 tpg|BK006945.2| 205583 + tpg|BK006945.2| 205943 - INS 
 tpg|BK006945.2| 202313 + tpg|BK006945.2| 202154 - INS 
 tpg|BK006936.2| 517425 + tpg|BK006936.2| 516923 - INS 
 tpg|BK006936.2| 603054 + tpg|BK006936.2| 602907 - INS 
 tpg|BK006936.2| 383156 + tpg|BK006936.2| 382697 - INS 
 tpg|BK006945.2| 116030 + tpg|BK006945.2| 116556 - INS 
 tpg|BK006936.2| 228997 + tpg|BK006936.2| 228589 - INS 
 tpg|BK006945.2| 363039 + tpg|BK006945.2| 362907 - INS 
 tpg|BK006936.2| 533203 + tpg|BK006936.2| 533392 - INS 
 tpg|BK006936.2| 430828 + tpg|BK006936.2| 430587 - INS 
 tpg|BK006936.2| 422012 + tpg|BK006936.2| 421644 - INS 
 tpg|BK006945.2| 198690 + tpg|BK006945.2| 198035 - INS 
 tpg|BK006936.2| 537961 + tpg|BK006936.2| 537614 - INS 
 tpg|BK006936.2| 792858 + tpg|BK006936.2| 792258 - INS 
 tpg|BK006936.2| 445727 + tpg|BK006936.2| 445532 - INS 
 tpg|BK006936.2| 47186 + tpg|BK006936.2| 46594 - INS 
 tpg|BK006936.2| 453359 + tpg|BK006936.2| 453383 - INS 
 tpg|BK006936.2| 418033 + tpg|BK006936.2| 417724 - INS 
 tpg|BK006936.2| 768066 + tpg|BK006936.2| 767567 - INS 
 tpg|BK006936.2| 62187 + tpg|BK006936.2| 61580 - INS 
 tpg|BK006945.2| 527802 + tpg|BK006945.2| 527117 - INS 
 tpg|BK006936.2| 398906 + tpg|BK006936.2| 399335 - INS 
 tpg|BK006945.2| 298382 + tpg|BK006945.2| 298022 - INS 
 tpg|BK006936.2| 66812 + tpg|BK006936.2| 67553 - INS 
 tpg|BK006936.2| 61633 + tpg|BK006936.2| 60922 - INS 
 tpg|BK006945.2| 1033021 + tpg|BK006945.2| 1033075 - INS 
 tpg|BK006936.2| 52745 + tpg|BK006936.2| 52538 - INS 
 tpg|BK006945.2| 890400 + tpg|BK006945.2| 890179 - INS 
 tpg|BK006936.2| 113991 + tpg|BK006936.2| 113817 - INS 
 tpg|BK006936.2| 716546 + tpg|BK006936.2| 715998 - INS 
 tpg|BK006936.2| 363780 + tpg|BK006936.2| 363595 - INS 
 tpg|BK006945.2| 170449 + tpg|BK006945.2| 170401 - INS 
 tpg|BK006936.2| 96528 + tpg|BK006936.2| 96520 - INS 
 tpg|BK006945.2| 710119 + tpg|BK006945.2| 709672 - INS 
 tpg|BK006936.2| 54232 + tpg|BK006936.2| 53644 - INS 
 tpg|BK006936.2| 162680 + tpg|BK006936.2| 162983 - INS 
 tpg|BK006936.2| 79580 + tpg|BK006936.2| 79580 - INS 
 tpg|BK006936.2| 446996 + tpg|BK006936.2| 446823 - INS 
 tpg|BK006945.2| 759518 + tpg|BK006945.2| 759391 - INS 
 tpg|BK006936.2| 697142 + tpg|BK006936.2| 696516 - INS 
 tpg|BK006936.2| 196517 + tpg|BK006936.2| 196387 - INS 
 tpg|BK006936.2| 766305 + tpg|BK006936.2| 766670 - INS 
 tpg|BK006945.2| 765259 + tpg|BK006945.2| 764915 - INS 
 tpg|BK006936.2| 586363 + tpg|BK006936.2| 585692 - INS 
 tpg|BK006936.2| 128599 + tpg|BK006936.2| 128456 - INS 
 tpg|BK006945.2| 613791 + tpg|BK006945.2| 613051 - INS 
 tpg|BK006936.2| 323937 + tpg|BK006936.2| 323977 - INS 
 tpg|BK006936.2| 140730 + tpg|BK006936.2| 140425 - INS 
 tpg|BK006945.2| 303491 + tpg|BK006945.2| 303835 - INS 
 tpg|BK006936.2| 75633 + tpg|BK006936.2| 74908 - INS 
 tpg|BK006945.2| 141049 + tpg|BK006945.2| 140339 - INS 
 tpg|BK006945.2| 632502 + tpg|BK006945.2| 632212 - INS 
 tpg|BK006936.2| 540489 + tpg|BK006936.2| 540550 - INS 
 tpg|BK006936.2| 469161 + tpg|BK006936.2| 468734 - INS 
 tpg|BK006936.2| 298395 + tpg|BK006936.2| 297990 - INS 
 tpg|BK006945.2| 810799 + tpg|BK006945.2| 810631 - INS 
 tpg|BK006945.2| 500327 + tpg|BK006945.2| 500292 - INS 
 tpg|BK006936.2| 469724 + tpg|BK006936.2| 469411 - INS 
 tpg|BK006936.2| 461638 + tpg|BK006936.2| 461401 - INS 
 tpg|BK006945.2| 315437 + tpg|BK006945.2| 316057 - INS 
 tpg|BK006936.2| 695534 + tpg|BK006936.2| 694900 - INS 
 tpg|BK006936.2| 289398 + tpg|BK006936.2| 289110 - INS 
 tpg|BK006945.2| 823792 + tpg|BK006945.2| 823714 - INS 
 tpg|BK006936.2| 688187 + tpg|BK006936.2| 688070 - INS 
 tpg|BK006936.2| 169020 + tpg|BK006936.2| 169372 - INS 
 tpg|BK006936.2| 220083 + tpg|BK006936.2| 219746 - INS 
 tpg|BK006945.2| 791000 + tpg|BK006945.2| 791211 - INS 
 tpg|BK006936.2| 216380 + tpg|BK006936.2| 216148 - INS 
 tpg|BK006945.2| 16222 + tpg|BK006945.2| 15819 - INS 
 tpg|BK006936.2| 762849 + tpg|BK006936.2| 763170 - INS 
 tpg|BK006945.2| 803330 + tpg|BK006945.2| 803162 - INS 
 tpg|BK006936.2| 443879 + tpg|BK006936.2| 443746 - INS 
 tpg|BK006945.2| 264388 + tpg|BK006945.2| 264070 - INS 
 tpg|BK006945.2| 286640 + tpg|BK006945.2| 286709 - INS 
 tpg|BK006945.2| 113285 + tpg|BK006945.2| 112537 - INS 
 tpg|BK006945.2| 548746 + tpg|BK006945.2| 548550 - INS 
 tpg|BK006936.2| 637774 + tpg|BK006936.2| 637406 - INS 
 tpg|BK006936.2| 413126 + tpg|BK006936.2| 412711 - INS 
 tpg|BK006945.2| 586640 + tpg|BK006945.2| 586512 - INS 
 tpg|BK006936.2| 532525 + tpg|BK006936.2| 532406 - INS 
 tpg|BK006945.2| 271132 + tpg|BK006945.2| 271829 - INS 
 tpg|BK006936.2| 416108 + tpg|BK006936.2| 415526 - INS 
 tpg|BK006936.2| 782513 + tpg|BK006936.2| 782827 - INS 
 tpg|BK006936.2| 179876 + tpg|BK006936.2| 179407 - INS 
 tpg|BK006945.2| 574128 + tpg|BK006945.2| 573838 - INS 
 tpg|BK006936.2| 683620 + tpg|BK006936.2| 683306 - INS 
 tpg|BK006945.2| 663812 + tpg|BK006945.2| 664257 - INS 
 tpg|BK006936.2| 525327 + tpg|BK006936.2| 525507 - INS 
 tpg|BK006936.2| 39883 + tpg|BK006936.2| 39601 - INS 
 tpg|BK006936.2| 111087 + tpg|BK006936.2| 110759 - INS 
 tpg|BK006936.2| 290351 + tpg|BK006936.2| 290310 - INS 
 tpg|BK006936.2| 575199 + tpg|BK006936.2| 575290 - INS 
 tpg|BK006936.2| 284003 + tpg|BK006936.2| 283803 - INS 
 tpg|BK006936.2| 321444 + tpg|BK006936.2| 321093 - INS 
 tpg|BK006945.2| 448528 + tpg|BK006945.2| 448774 - INS 
 tpg|BK006936.2| 89874 + tpg|BK006936.2| 90062 - INS 
 tpg|BK006936.2| 805636 + tpg|BK006936.2| 805087 - INS 
 tpg|BK006945.2| 717995 + tpg|BK006945.2| 718247 - INS 
 tpg|BK006936.2| 129377 + tpg|BK006936.2| 129824 - INS 
 tpg|BK006936.2| 279769 + tpg|BK006936.2| 279386 - INS 
 tpg|BK006936.2| 92749 + tpg|BK006936.2| 92104 - INS 
 tpg|BK006936.2| 654963 + tpg|BK006936.2| 655182 - INS 
 tpg|BK006936.2| 545396 + tpg|BK006936.2| 545616 - INS 
 tpg|BK006936.2| 29598 + tpg|BK006936.2| 29419 - INS 
 tpg|BK006936.2| 245953 + tpg|BK006936.2| 245780 - INS 
 tpg|BK006945.2| 114254 + tpg|BK006945.2| 113999 - INS 
 tpg|BK006936.2| 402605 + tpg|BK006936.2| 401893 - INS 
 tpg|BK006936.2| 429926 + tpg|BK006936.2| 429668 - INS 
 tpg|BK006936.2| 9546 + tpg|BK006936.2| 9691 - INS 
 tpg|BK006936.2| 521551 + tpg|BK006936.2| 521017 - INS 
 tpg|BK006945.2| 850541 + tpg|BK006945.2| 850380 - INS 
 tpg|BK006936.2| 586822 + tpg|BK006936.2| 586595 - INS 
 tpg|BK006936.2| 38136 + tpg|BK006936.2| 37953 - INS 
 tpg|BK006936.2| 124357 + tpg|BK006936.2| 124051 - INS GAAA
 tpg|BK006936.2| 301343 + tpg|BK006936.2| 301253 - INS 
 tpg|BK006945.2| 634721 + tpg|BK006945.2| 634502 - INS 
 tpg|BK006936.2| 436621 + tpg|BK006936.2| 436091 - INS 
 tpg|BK006936.2| 636004 + tpg|BK006936.2| 635759 - INS 
 tpg|BK006945.2| 579730 + tpg|BK006945.2| 579215 - INS 
 tpg|BK006936.2| 155772 + tpg|BK006936.2| 155717 - INS 
 tpg|BK006936.2| 188910 + tpg|BK006936.2| 188785 - INS 
 tpg|BK006936.2| 8663 + tpg|BK006936.2| 8321 - INS 
 tpg|BK006936.2| 507144 + tpg|BK006936.2| 507068 - INS 
 tpg|BK006945.2| 692863 + tpg|BK006945.2| 692386 - INS 
 tpg|BK006945.2| 1008294 + tpg|BK006945.2| 1008978 - INS 
 tpg|BK006945.2| 846414 + tpg|BK006945.2| 846730 - INS 
 tpg|BK006945.2| 675699 + tpg|BK006945.2| 675363 - INS 
 tpg|BK006945.2| 966274 + tpg|BK006945.2| 967010 - INS 
 tpg|BK006945.2| 668368 + tpg|BK006945.2| 669086 - INS 
 tpg|BK006945.2| 920603 + tpg|BK006945.2| 919923 - INS 
 tpg|BK006945.2| 184271 + tpg|BK006945.2| 184904 - INS 
 tpg|BK006945.2| 200962 + tpg|BK006945.2| 200583 - INS 
 tpg|BK006945.2| 862364 + tpg|BK006945.2| 861940 - INS 
 tpg|BK006945.2| 290003 + tpg|BK006945.2| 289853 - INS 
 tpg|BK006945.2| 697017 + tpg|BK006945.2| 696571 - INS 
 tpg|BK006945.2| 899704 + tpg|BK006945.2| 899189 - INS 
 tpg|BK006945.2| 172653 + tpg|BK006945.2| 172196 - INS 
 tpg|BK006945.2| 40826 + tpg|BK006945.2| 40262 - INS 
 tpg|BK006945.2| 1029671 + tpg|BK006945.2| 1029009 - INS 
 tpg|BK006945.2| 931990 + tpg|BK006945.2| 932027 - INS 
 tpg|BK006945.2| 1023153 + tpg|BK006945.2| 1023058 - INS 
 tpg|BK006945.2| 62882 + tpg|BK006945.2| 62549 - INS 
 tpg|BK006945.2| 764565 + tpg|BK006945.2| 763923 - INS 
 tpg|BK006945.2| 775687 + tpg|BK006945.2| 776395 - INS 
 tpg|BK006945.2| 310556 + tpg|BK006945.2| 309906 - INS 
 tpg|BK006945.2| 624166 + tpg|BK006945.2| 623614 - INS 
 tpg|BK006945.2| 954121 + tpg|BK006945.2| 954416 - INS 
 tpg|BK006945.2| 822282 + tpg|BK006945.2| 822830 - INS 
 tpg|BK006945.2| 17553 + tpg|BK006945.2| 17178 - INS 
 tpg|BK006945.2| 590256 + tpg|BK006945.2| 590597 - INS 
 tpg|BK006945.2| 77306 + tpg|BK006945.2| 76711 - INS 
 tpg|BK006945.2| 549546 + tpg|BK006945.2| 549737 - INS 
 tpg|BK006945.2| 551762 + tpg|BK006945.2| 551612 - INS 
 tpg|BK006945.2| 585069 + tpg|BK006945.2| 585691 - INS 
 tpg|BK006945.2| 531925 + tpg|BK006945.2| 532191 - INS GCTTGCA
 tpg|BK006945.2| 814247 + tpg|BK006945.2| 814509 - INS AAT
 tpg|BK006944.2| 6808 + tpg|BK006944.2| 6424 - INS 
 tpg|BK006945.2| 805706 + tpg|BK006945.2| 805671 - INS 
 tpg|BK006945.2| 800656 + tpg|BK006945.2| 800941 - INS 
 tpg|BK006945.2| 299664 + tpg|BK006945.2| 299686 - INS 
 tpg|BK006945.2| 233593 + tpg|BK006945.2| 233625 - INS 
 tpg|BK006944.2| 572216 + tpg|BK006944.2| 572903 - INS 
 tpg|BK006945.2| 506421 + tpg|BK006945.2| 506326 - INS 
 tpg|BK006945.2| 859571 + tpg|BK006945.2| 859467 - INS 
 tpg|BK006944.2| 87459 + tpg|BK006944.2| 87723 - INS 
 tpg|BK006945.2| 639877 + tpg|BK006945.2| 639425 - INS 
 tpg|BK006945.2| 149887 + tpg|BK006945.2| 149368 - INS 
 tpg|BK006945.2| 748732 + tpg|BK006945.2| 748852 - INS 
 tpg|BK006944.2| 528843 + tpg|BK006944.2| 529065 - INS 
 tpg|BK006945.2| 647214 + tpg|BK006945.2| 647212 - INS 
 tpg|BK006944.2| 519635 + tpg|BK006944.2| 519840 - INS 
 tpg|BK006945.2| 728597 + tpg|BK006945.2| 728870 - INS 
 tpg|BK006945.2| 155443 + tpg|BK006945.2| 155199 - INS 
 tpg|BK006944.2| 485918 + tpg|BK006944.2| 486479 - INS 
 tpg|BK006945.2| 1021670 + tpg|BK006945.2| 1021351 - INS 
 tpg|BK006944.2| 171199 + tpg|BK006944.2| 170930 - INS 
 tpg|BK006945.2| 1033891 + tpg|BK006945.2| 1034397 - INS 
 tpg|BK006945.2| 687947 + tpg|BK006945.2| 687356 - INS 
 tpg|BK006945.2| 910098 + tpg|BK006945.2| 909738 - INS 
 tpg|BK006945.2| 721528 + tpg|BK006945.2| 721352 - INS 
 tpg|BK006944.2| 58975 + tpg|BK006944.2| 59148 - INS 
 tpg|BK006945.2| 956521 + tpg|BK006945.2| 956449 - INS 
 tpg|BK006945.2| 57757 + tpg|BK006945.2| 58330 - INS 
 tpg|BK006944.2| 367015 + tpg|BK006944.2| 366850 - INS 
 tpg|BK006945.2| 526791 + tpg|BK006945.2| 526602 - INS 
 tpg|BK006944.2| 286157 + tpg|BK006944.2| 286236 - INS 
 tpg|BK006945.2| 71578 + tpg|BK006945.2| 70828 - INS 
 tpg|BK006944.2| 93789 + tpg|BK006944.2| 93130 - INS 
 tpg|BK006945.2| 864704 + tpg|BK006945.2| 864076 - INS 
 tpg|BK006945.2| 567112 + tpg|BK006945.2| 566928 - INS 
 tpg|BK006945.2| 905478 + tpg|BK006945.2| 905102 - INS 
 tpg|BK006944.2| 230253 + tpg|BK006944.2| 230346 - INS 
 tpg|BK006944.2| 116049 + tpg|BK006944.2| 115655 - INS 
 tpg|BK006945.2| 284760 + tpg|BK006945.2| 284674 - INS 
 tpg|BK006944.2| 322942 + tpg|BK006944.2| 322455 - INS 
 tpg|BK006945.2| 987521 + tpg|BK006945.2| 987176 - INS 
 tpg|BK006949.2| 763242 + tpg|BK006949.2| 763231 - INS 
 tpg|BK006944.2| 59810 + tpg|BK006944.2| 60458 - INS 
 tpg|BK006945.2| 985152 + tpg|BK006945.2| 984955 - INS 
 tpg|BK006945.2| 964583 + tpg|BK006945.2| 964336 - INS 
 tpg|BK006945.2| 134314 + tpg|BK006945.2| 134818 - INS 
 tpg|BK006945.2| 123420 + tpg|BK006945.2| 123315 - INS 
 tpg|BK006949.2| 392628 + tpg|BK006949.2| 393111 - INS 
 tpg|BK006945.2| 941173 + tpg|BK006945.2| 940876 - INS 
 tpg|BK006944.2| 594903 + tpg|BK006944.2| 594316 - INS 
 tpg|BK006945.2| 919138 + tpg|BK006945.2| 918523 - INS 
 tpg|BK006945.2| 383902 + tpg|BK006945.2| 383266 - INS 
 tpg|BK006945.2| 378711 + tpg|BK006945.2| 379046 - INS 
 tpg|BK006949.2| 402951 + tpg|BK006949.2| 402812 - INS 
 tpg|BK006944.2| 16857 + tpg|BK006944.2| 16455 - INS 
 tpg|BK006945.2| 1042288 + tpg|BK006945.2| 1042272 - INS 
 tpg|BK006945.2| 226009 + tpg|BK006945.2| 225238 - INS 
 tpg|BK006944.2| 356654 + tpg|BK006944.2| 357221 - INS 
 tpg|BK006945.2| 45111 + tpg|BK006945.2| 44372 - INS 
 tpg|BK006944.2| 362313 + tpg|BK006944.2| 361926 - INS 
 tpg|BK006945.2| 891226 + tpg|BK006945.2| 891433 - INS 
 tpg|BK006944.2| 73955 + tpg|BK006944.2| 73225 - INS 
 tpg|BK006945.2| 194154 + tpg|BK006945.2| 194595 - INS 
 tpg|BK006945.2| 183627 + tpg|BK006945.2| 183237 - INS 
 tpg|BK006944.2| 149645 + tpg|BK006944.2| 149149 - INS 
 tpg|BK006945.2| 991391 + tpg|BK006945.2| 991341 - INS 
 tpg|BK006944.2| 477136 + tpg|BK006944.2| 477596 - INS 
 tpg|BK006945.2| 182865 + tpg|BK006945.2| 182481 - INS 
 tpg|BK006945.2| 247813 + tpg|BK006945.2| 247908 - INS 
 tpg|BK006944.2| 479954 + tpg|BK006944.2| 479866 - INS 
 tpg|BK006945.2| 296868 + tpg|BK006945.2| 296138 - INS 
 tpg|BK006945.2| 177587 + tpg|BK006945.2| 177415 - INS 
 tpg|BK006945.2| 358279 + tpg|BK006945.2| 357860 - INS 
 tpg|BK006944.2| 617003 + tpg|BK006944.2| 616354 - INS 
 tpg|BK006945.2| 212702 + tpg|BK006945.2| 213465 - INS 
 tpg|BK006945.2| 146036 + tpg|BK006945.2| 145393 - INS 
 tpg|BK006944.2| 499031 + tpg|BK006944.2| 498333 - INS 
 tpg|BK006945.2| 1046035 + tpg|BK006945.2| 1045593 - INS 
 tpg|BK006945.2| 497680 + tpg|BK006945.2| 498143 - INS 
 tpg|BK006944.2| 496596 + tpg|BK006944.2| 495922 - INS 
 tpg|BK006945.2| 769090 + tpg|BK006945.2| 769827 - INS 
 tpg|BK006944.2| 518362 + tpg|BK006944.2| 518567 - INS 
 tpg|BK006945.2| 509109 + tpg|BK006945.2| 508816 - INS 
 tpg|BK006945.2| 784517 + tpg|BK006945.2| 784444 - INS 
 tpg|BK006945.2| 535789 + tpg|BK006945.2| 535166 - INS 
 tpg|BK006949.2| 343225 + tpg|BK006949.2| 342937 - INS 
 tpg|BK006945.2| 66212 + tpg|BK006945.2| 65968 - INS 
 tpg|BK006945.2| 968854 + tpg|BK006945.2| 968271 - INS 
 tpg|BK006945.2| 845027 + tpg|BK006945.2| 844265 - INS 
 tpg|BK006945.2| 554729 + tpg|BK006945.2| 554306 - INS 
 tpg|BK006945.2| 660578 + tpg|BK006945.2| 660299 - INS 
 tpg|BK006944.2| 453709 + tpg|BK006944.2| 453161 - INS 
 tpg|BK006945.2| 808808 + tpg|BK006945.2| 808244 - INS 
 tpg|BK006949.2| 791079 + tpg|BK006949.2| 790430 - INS 
 tpg|BK006944.2| 448889 + tpg|BK006944.2| 448896 - INS 
 tpg|BK006945.2| 602708 + tpg|BK006945.2| 602502 - INS 
 tpg|BK006945.2| 91248 + tpg|BK006945.2| 90509 - INS 
 tpg|BK006949.2| 465931 + tpg|BK006949.2| 465663 - INS 
 tpg|BK006945.2| 965764 + tpg|BK006945.2| 965401 - INS 
 tpg|BK006944.2| 562403 + tpg|BK006944.2| 562012 - INS 
 tpg|BK006945.2| 995631 + tpg|BK006945.2| 995513 - INS 
 tpg|BK006949.2| 553486 + tpg|BK006949.2| 553149 - INS 
 tpg|BK006945.2| 359269 + tpg|BK006945.2| 359365 - INS 
 tpg|BK006949.2| 76737 + tpg|BK006949.2| 76321 - INS 
 tpg|BK006945.2| 1062976 + tpg|BK006945.2| 1062323 - INS 
 tpg|BK006945.2| 251739 + tpg|BK006945.2| 251193 - INS 
 tpg|BK006944.2| 608820 + tpg|BK006944.2| 608372 - INS 
 tpg|BK006945.2| 1061564 + tpg|BK006945.2| 1061215 - INS 
 tpg|BK006949.2| 194288 + tpg|BK006949.2| 194110 - INS 
 tpg|BK006945.2| 915408 + tpg|BK006945.2| 915214 - INS 
 tpg|BK006945.2| 565056 + tpg|BK006945.2| 565137 - INS 
 tpg|BK006944.2| 240292 + tpg|BK006944.2| 239894 - INS 
 tpg|BK006945.2| 1058814 + tpg|BK006945.2| 1058786 - INS 
 tpg|BK006949.2| 753973 + tpg|BK006949.2| 753231 - INS 
 tpg|BK006945.2| 583052 + tpg|BK006945.2| 582880 - INS 
 tpg|BK006945.2| 557447 + tpg|BK006945.2| 557426 - INS 
 tpg|BK006945.2| 42227 + tpg|BK006945.2| 42888 - INS 
 tpg|BK006944.2| 317392 + tpg|BK006944.2| 317088 - INS 
 tpg|BK006949.2| 827440 + tpg|BK006949.2| 827131 - INS 
 tpg|BK006945.2| 55627 + tpg|BK006945.2| 55101 - INS 
 tpg|BK006944.2| 14970 + tpg|BK006944.2| 14338 - INS 
 tpg|BK006945.2| 609567 + tpg|BK006945.2| 609252 - INS 
 tpg|BK006945.2| 924033 + tpg|BK006945.2| 924170 - INS 
 tpg|BK006944.2| 525006 + tpg|BK006944.2| 524836 - INS 
 tpg|BK006945.2| 675216 + tpg|BK006945.2| 674700 - INS 
 tpg|BK006945.2| 108969 + tpg|BK006945.2| 109445 - INS 
 tpg|BK006945.2| 444110 + tpg|BK006945.2| 444533 - INS 
 tpg|BK006944.2| 457268 + tpg|BK006944.2| 457543 - INS 
 tpg|BK006945.2| 244581 + tpg|BK006945.2| 243881 - INS 
 tpg|BK006945.2| 428102 + tpg|BK006945.2| 427584 - INS 
 tpg|BK006949.2| 680448 + tpg|BK006949.2| 680138 - INS 
 tpg|BK006945.2| 925219 + tpg|BK006945.2| 924924 - INS 
 tpg|BK006944.2| 435517 + tpg|BK006944.2| 435162 - INS 
 tpg|BK006945.2| 345040 + tpg|BK006945.2| 345282 - INS 
 tpg|BK006945.2| 285568 + tpg|BK006945.2| 286311 - INS 
 tpg|BK006944.2| 239500 + tpg|BK006944.2| 239176 - INS 
 tpg|BK006949.2| 501734 + tpg|BK006949.2| 502464 - INS 
 tpg|BK006944.2| 464732 + tpg|BK006944.2| 464612 - INS 
 tpg|BK006945.2| 1019094 + tpg|BK006945.2| 1019832 - INS 
 tpg|BK006945.2| 334710 + tpg|BK006945.2| 334093 - INS 
 tpg|BK006944.2| 619464 + tpg|BK006944.2| 619308 - INS 
 tpg|BK006949.2| 75995 + tpg|BK006949.2| 75511 - INS 
 tpg|BK006945.2| 193133 + tpg|BK006945.2| 193344 - INS 
 tpg|BK006945.2| 740114 + tpg|BK006945.2| 740167 - INS 
 tpg|BK006944.2| 168701 + tpg|BK006944.2| 168304 - INS 
 tpg|BK006945.2| 343535 + tpg|BK006945.2| 343843 - INS 
 tpg|BK006949.2| 511860 + tpg|BK006949.2| 512263 - INS 
 tpg|BK006944.2| 319447 + tpg|BK006944.2| 318722 - INS 
 tpg|BK006945.2| 1027449 + tpg|BK006945.2| 1027020 - INS 
 tpg|BK006945.2| 348716 + tpg|BK006945.2| 349009 - INS 
 tpg|BK006945.2| 31056 + tpg|BK006945.2| 30805 - INS 
 tpg|BK006945.2| 268526 + tpg|BK006945.2| 268478 - INS 
 tpg|BK006944.2| 586215 + tpg|BK006944.2| 585441 - INS 
 tpg|BK006949.2| 184674 + tpg|BK006949.2| 185250 - INS 
 tpg|BK006945.2| 300487 + tpg|BK006945.2| 300974 - INS 
 tpg|BK006944.2| 646576 + tpg|BK006944.2| 647231 - INS 
 tpg|BK006945.2| 305975 + tpg|BK006945.2| 305638 - INS 
 tpg|BK006949.2| 628366 + tpg|BK006949.2| 628685 - INS 
 tpg|BK006945.2| 308566 + tpg|BK006945.2| 308450 - INS 
 tpg|BK006944.2| 531540 + tpg|BK006944.2| 532000 - INS 
 tpg|BK006945.2| 406555 + tpg|BK006945.2| 405837 - INS 
 tpg|BK006945.2| 405830 + tpg|BK006945.2| 405364 - INS 
 tpg|BK006944.2| 558595 + tpg|BK006944.2| 557951 - INS 
 tpg|BK006949.2| 518228 + tpg|BK006949.2| 518368 - INS 
 tpg|BK006944.2| 440974 + tpg|BK006944.2| 440885 - INS 
 tpg|BK006945.2| 439595 + tpg|BK006945.2| 440249 - INS 
 tpg|BK006945.2| 51435 + tpg|BK006945.2| 51060 - INS 
 tpg|BK006949.2| 289436 + tpg|BK006949.2| 289249 - INS 
 tpg|BK006944.2| 570746 + tpg|BK006944.2| 570511 - INS 
 tpg|BK006945.2| 701255 + tpg|BK006945.2| 700775 - INS 
 tpg|BK006949.2| 161444 + tpg|BK006949.2| 160839 - INS 
 tpg|BK006945.2| 513512 + tpg|BK006945.2| 513375 - INS 
 tpg|BK006944.2| 37490 + tpg|BK006944.2| 37743 - INS 
 tpg|BK006945.2| 85107 + tpg|BK006945.2| 84815 - INS 
 tpg|BK006944.2| 476015 + tpg|BK006944.2| 475661 - INS 
 tpg|BK006944.2| 30794 + tpg|BK006944.2| 31473 - INS 
 tpg|BK006945.2| 63996 + tpg|BK006945.2| 63500 - INS 
 tpg|BK006945.2| 686554 + tpg|BK006945.2| 686348 - INS 
 tpg|BK006945.2| 555546 + tpg|BK006945.2| 555312 - INS 
 tpg|BK006949.2| 359083 + tpg|BK006949.2| 358586 - INS 
 tpg|BK006945.2| 307471 + tpg|BK006945.2| 307403 - INS 
 tpg|BK006945.2| 900145 + tpg|BK006945.2| 900550 - INS 
 tpg|BK006944.2| 379992 + tpg|BK006944.2| 380014 - INS 
 tpg|BK006945.2| 910856 + tpg|BK006945.2| 910404 - INS 
 tpg|BK006945.2| 914869 + tpg|BK006945.2| 914394 - INS 
 tpg|BK006945.2| 409032 + tpg|BK006945.2| 409215 - INS 
 tpg|BK006944.2| 488158 + tpg|BK006944.2| 488081 - INS 
 tpg|BK006949.2| 228132 + tpg|BK006949.2| 227448 - INS 
 tpg|BK006945.2| 162252 + tpg|BK006945.2| 161830 - INS 
 tpg|BK006945.2| 883210 + tpg|BK006945.2| 882930 - INS 
 tpg|BK006949.2| 835159 + tpg|BK006949.2| 835227 - INS 
 tpg|BK006944.2| 351216 + tpg|BK006944.2| 350543 - INS 
 tpg|BK006945.2| 1043093 + tpg|BK006945.2| 1043078 - INS 
 tpg|BK006945.2| 667897 + tpg|BK006945.2| 668420 - INS 
 tpg|BK006949.2| 738433 + tpg|BK006949.2| 738608 - INS 
 tpg|BK006945.2| 722340 + tpg|BK006945.2| 721757 - INS 
 tpg|BK006944.2| 369979 + tpg|BK006944.2| 369529 - INS 
 tpg|BK006945.2| 335330 + tpg|BK006945.2| 334688 - INS 
 tpg|BK006945.2| 755392 + tpg|BK006945.2| 755102 - INS 
 tpg|BK006944.2| 340612 + tpg|BK006944.2| 340408 - INS 
 tpg|BK006944.2| 101051 + tpg|BK006944.2| 100749 - INS 
 tpg|BK006949.2| 677105 + tpg|BK006949.2| 677657 - INS 
 tpg|BK006945.2| 32788 + tpg|BK006945.2| 32582 - INS 
 tpg|BK006945.2| 492925 + tpg|BK006945.2| 492230 - INS 
 tpg|BK006945.2| 493485 + tpg|BK006945.2| 492748 - INS 
 tpg|BK006949.2| 31859 + tpg|BK006949.2| 31301 - INS 
 tpg|BK006945.2| 950852 + tpg|BK006945.2| 950354 - INS 
 tpg|BK006945.2| 1053809 + tpg|BK006945.2| 1053483 - INS 
 tpg|BK006944.2| 655853 + tpg|BK006944.2| 656281 - INS 
 tpg|BK006949.2| 199435 + tpg|BK006949.2| 198733 - INS 
 tpg|BK006945.2| 892531 + tpg|BK006945.2| 892017 - INS 
 tpg|BK006945.2| 238069 + tpg|BK006945.2| 237870 - INS 
 tpg|BK006945.2| 614998 + tpg|BK006945.2| 614619 - INS 
 tpg|BK006944.2| 600654 + tpg|BK006944.2| 601150 - INS 
 tpg|BK006945.2| 852744 + tpg|BK006945.2| 852258 - INS 
 tpg|BK006949.2| 68797 + tpg|BK006949.2| 68577 - INS 
 tpg|BK006945.2| 770665 + tpg|BK006945.2| 771028 - INS 
 tpg|BK006944.2| 328271 + tpg|BK006944.2| 328917 - INS ACT
 tpg|BK006945.2| 848679 + tpg|BK006945.2| 848368 - INS 
 tpg|BK006949.2| 921367 + tpg|BK006949.2| 921155 - INS 
 tpg|BK006945.2| 108404 + tpg|BK006945.2| 108388 - INS 
 tpg|BK006949.2| 197913 + tpg|BK006949.2| 198057 - INS 
 tpg|BK006944.2| 194048 + tpg|BK006944.2| 193355 - INS 
 tpg|BK006945.2| 926732 + tpg|BK006945.2| 927338 - INS 
 tpg|BK006944.2| 21843 + tpg|BK006944.2| 21177 - INS 
 tpg|BK006945.2| 1056924 + tpg|BK006945.2| 1056784 - INS 
 tpg|BK006949.2| 188693 + tpg|BK006949.2| 188036 - INS 
 tpg|BK006945.2| 1050887 + tpg|BK006945.2| 1050461 - INS 
 tpg|BK006944.2| 247599 + tpg|BK006944.2| 247018 - INS 
 tpg|BK006945.2| 317224 + tpg|BK006945.2| 317720 - INS 
 tpg|BK006945.2| 27409 + tpg|BK006945.2| 27083 - INS 
 tpg|BK006944.2| 535536 + tpg|BK006944.2| 535431 - INS 
 tpg|BK006945.2| 1030387 + tpg|BK006945.2| 1029819 - INS 
 tpg|BK006949.2| 82223 + tpg|BK006949.2| 81520 - INS 
 tpg|BK006944.2| 345556 + tpg|BK006944.2| 345039 - INS 
 tpg|BK006945.2| 857895 + tpg|BK006945.2| 857545 - INS 
 tpg|BK006944.2| 122408 + tpg|BK006944.2| 122500 - INS 
 tpg|BK006945.2| 948351 + tpg|BK006945.2| 947783 - INS 
 tpg|BK006945.2| 666485 + tpg|BK006945.2| 666258 - INS 
 tpg|BK006949.2| 158379 + tpg|BK006949.2| 158345 - INS 
 tpg|BK006944.2| 63544 + tpg|BK006944.2| 64040 - INS 
 tpg|BK006945.2| 173925 + tpg|BK006945.2| 173853 - INS 
 tpg|BK006949.2| 407109 + tpg|BK006949.2| 406776 - INS 
 tpg|BK006945.2| 906684 + tpg|BK006945.2| 906433 - INS 
 tpg|BK006945.2| 738218 + tpg|BK006945.2| 737817 - INS 
 tpg|BK006949.2| 455556 + tpg|BK006949.2| 455207 - INS 
 tpg|BK006945.2| 187593 + tpg|BK006945.2| 186946 - INS 
 tpg|BK006945.2| 209126 + tpg|BK006945.2| 209645 - INS 
 tpg|BK006944.2| 463287 + tpg|BK006944.2| 463266 - INS 
 tpg|BK006945.2| 868985 + tpg|BK006945.2| 868416 - INS 
 tpg|BK006945.2| 836273 + tpg|BK006945.2| 836244 - INS 
 tpg|BK006945.2| 178540 + tpg|BK006945.2| 177987 - INS 
 tpg|BK006944.2| 383708 + tpg|BK006944.2| 383466 - INS 
 tpg|BK006949.2| 360749 + tpg|BK006949.2| 360749 - INS 
 tpg|BK006944.2| 246557 + tpg|BK006944.2| 246082 - INS 
 tpg|BK006945.2| 83203 + tpg|BK006945.2| 83115 - INS 
 tpg|BK006945.2| 546117 + tpg|BK006945.2| 545524 - INS 
 tpg|BK006945.2| 902187 + tpg|BK006945.2| 902063 - INS 
 tpg|BK006944.2| 474406 + tpg|BK006944.2| 474365 - INS 
 tpg|BK006949.2| 609717 + tpg|BK006949.2| 609356 - INS 
 tpg|BK006945.2| 813612 + tpg|BK006945.2| 812926 - INS 
 tpg|BK006949.2| 786494 + tpg|BK006949.2| 786911 - INS 
 tpg|BK006944.2| 282780 + tpg|BK006944.2| 283383 - INS 
 tpg|BK006945.2| 809649 + tpg|BK006945.2| 809853 - INS 
 tpg|BK006944.2| 639886 + tpg|BK006944.2| 639993 - INS 
 tpg|BK006945.2| 624743 + tpg|BK006945.2| 624552 - INS 
 tpg|BK006949.2| 479604 + tpg|BK006949.2| 479067 - INS 
 tpg|BK006945.2| 115450 + tpg|BK006945.2| 115311 - INS 
 tpg|BK006945.2| 60784 + tpg|BK006945.2| 60869 - INS 
 tpg|BK006944.2| 17498 + tpg|BK006944.2| 17241 - INS 
 tpg|BK006945.2| 60080 + tpg|BK006945.2| 59865 - INS 
 tpg|BK006949.2| 686851 + tpg|BK006949.2| 687135 - INS 
 tpg|BK006945.2| 833679 + tpg|BK006945.2| 833459 - INS 
 tpg|BK006945.2| 842945 + tpg|BK006945.2| 842620 - INS 
 tpg|BK006945.2| 33640 + tpg|BK006945.2| 33710 - INS 
 tpg|BK006945.2| 661058 + tpg|BK006945.2| 661552 - INS 
 tpg|BK006945.2| 509692 + tpg|BK006945.2| 509880 - INS 
 tpg|BK006944.2| 423624 + tpg|BK006944.2| 423102 - INS 
 tpg|BK006945.2| 46504 + tpg|BK006945.2| 46426 - INS 
 tpg|BK006945.2| 936566 + tpg|BK006945.2| 936061 - INS 
 tpg|BK006945.2| 256513 + tpg|BK006945.2| 256062 - INS 
 tpg|BK006944.2| 494047 + tpg|BK006944.2| 494197 - INS 
 tpg|BK006945.2| 633124 + tpg|BK006945.2| 632917 - INS 
 tpg|BK006945.2| 407122 + tpg|BK006945.2| 407091 - INS 
 tpg|BK006944.2| 569376 + tpg|BK006944.2| 569377 - INS 
 tpg|BK006945.2| 324103 + tpg|BK006945.2| 323909 - INS 
 tpg|BK006945.2| 912267 + tpg|BK006945.2| 912363 - INS 
 tpg|BK006949.2| 447975 + tpg|BK006949.2| 447876 - INS 
 tpg|BK006945.2| 56792 + tpg|BK006945.2| 56482 - INS 
 tpg|BK006945.2| 433303 + tpg|BK006945.2| 433244 - INS 
 tpg|BK006945.2| 929287 + tpg|BK006945.2| 928743 - INS 
 tpg|BK006949.2| 863934 + tpg|BK006949.2| 863198 - INS 
 tpg|BK006945.2| 50844 + tpg|BK006945.2| 50152 - INS 
 tpg|BK006945.2| 717408 + tpg|BK006945.2| 717366 - INS 
 tpg|BK006945.2| 211044 + tpg|BK006945.2| 210293 - INS 
 tpg|BK006944.2| 513767 + tpg|BK006944.2| 513380 - INS 
 tpg|BK006945.2| 603598 + tpg|BK006945.2| 603124 - INS 
 tpg|BK006949.2| 187184 + tpg|BK006949.2| 187124 - INS 
 tpg|BK006945.2| 678148 + tpg|BK006945.2| 677842 - INS 
 tpg|BK006944.2| 95179 + tpg|BK006944.2| 95635 - INS 
 tpg|BK006945.2| 52661 + tpg|BK006945.2| 52234 - INS 
 tpg|BK006945.2| 1027845 + tpg|BK006945.2| 1027836 - INS 
 tpg|BK006945.2| 1026104 + tpg|BK006945.2| 1025828 - INS 
 tpg|BK006945.2| 994342 + tpg|BK006945.2| 993879 - INS 
 tpg|BK006944.2| 315332 + tpg|BK006944.2| 314641 - INS 
 tpg|BK006945.2| 546769 + tpg|BK006945.2| 546966 - INS 
 tpg|BK006945.2| 730530 + tpg|BK006945.2| 730809 - INS 
 tpg|BK006949.2| 821744 + tpg|BK006949.2| 821924 - INS 
 tpg|BK006944.2| 82247 + tpg|BK006944.2| 81524 - INS 
 tpg|BK006945.2| 708092 + tpg|BK006945.2| 707397 - INS 
 tpg|BK006945.2| 697967 + tpg|BK006945.2| 697390 - INS 
 tpg|BK006944.2| 288622 + tpg|BK006944.2| 288719 - INS 
 tpg|BK006949.2| 120580 + tpg|BK006949.2| 120499 - INS 
 tpg|BK006944.2| 404388 + tpg|BK006944.2| 403807 - INS 
 tpg|BK006944.2| 23603 + tpg|BK006944.2| 22922 - INS 
 tpg|BK006949.2| 319219 + tpg|BK006949.2| 319982 - INS 
 tpg|BK006949.2| 300669 + tpg|BK006949.2| 300664 - INS 
 tpg|BK006945.2| 883963 + tpg|BK006945.2| 884314 - INS 
 tpg|BK006944.2| 377919 + tpg|BK006944.2| 377215 - INS 
 tpg|BK006945.2| 865148 + tpg|BK006945.2| 865224 - INS 
 tpg|BK006944.2| 363768 + tpg|BK006944.2| 363096 - INS 
 tpg|BK006945.2| 752872 + tpg|BK006945.2| 752786 - INS 
 tpg|BK006945.2| 563378 + tpg|BK006945.2| 562696 - INS 
 tpg|BK006944.2| 203952 + tpg|BK006944.2| 203500 - INS 
 tpg|BK006945.2| 768088 + tpg|BK006945.2| 768135 - INS 
 tpg|BK006944.2| 272211 + tpg|BK006944.2| 272720 - INS 
 tpg|BK006945.2| 821119 + tpg|BK006945.2| 821822 - INS 
 tpg|BK006944.2| 384323 + tpg|BK006944.2| 384055 - INS 
 tpg|BK006945.2| 505785 + tpg|BK006945.2| 505328 - INS 
 tpg|BK006944.2| 251089 + tpg|BK006944.2| 251708 - INS 
 tpg|BK006945.2| 908792 + tpg|BK006945.2| 908698 - INS 
 tpg|BK006945.2| 438353 + tpg|BK006945.2| 438548 - INS 
 tpg|BK006945.2| 150634 + tpg|BK006945.2| 151011 - INS 
 tpg|BK006945.2| 740707 + tpg|BK006945.2| 741084 - INS 
 tpg|BK006944.2| 301651 + tpg|BK006944.2| 302220 - INS 
 tpg|BK006945.2| 658734 + tpg|BK006945.2| 658768 - INS 
 tpg|BK006945.2| 204860 + tpg|BK006945.2| 204444 - INS 
 tpg|BK006944.2| 134068 + tpg|BK006944.2| 134585 - INS 
 tpg|BK006945.2| 221180 + tpg|BK006945.2| 220865 - INS 
 tpg|BK006945.2| 911400 + tpg|BK006945.2| 911410 - INS 
 tpg|BK006949.2| 398403 + tpg|BK006949.2| 397630 - INS 
 tpg|BK006945.2| 5870 + tpg|BK006945.2| 5560 - INS 
 tpg|BK006944.2| 358031 + tpg|BK006944.2| 357982 - INS 
 tpg|BK006949.2| 373419 + tpg|BK006949.2| 373707 - INS 
 tpg|BK006944.2| 200313 + tpg|BK006944.2| 200137 - INS 
 tpg|BK006945.2| 263627 + tpg|BK006945.2| 263496 - INS 
 tpg|BK006944.2| 210974 + tpg|BK006944.2| 210217 - INS 
 tpg|BK006945.2| 153350 + tpg|BK006945.2| 153321 - INS 
 tpg|BK006945.2| 507352 + tpg|BK006945.2| 506993 - INS 
 tpg|BK006949.2| 73160 + tpg|BK006949.2| 73104 - INS 
 tpg|BK006944.2| 521494 + tpg|BK006944.2| 520997 - INS 
 tpg|BK006945.2| 961191 + tpg|BK006945.2| 961527 - INS 
 tpg|BK006945.2| 743067 + tpg|BK006945.2| 743542 - INS 
 tpg|BK006949.2| 497632 + tpg|BK006949.2| 498260 - INS 
 tpg|BK006945.2| 619139 + tpg|BK006945.2| 618790 - INS 
 tpg|BK006944.2| 314608 + tpg|BK006944.2| 313869 - INS 
 tpg|BK006945.2| 257119 + tpg|BK006945.2| 257295 - INS 
 tpg|BK006945.2| 614454 + tpg|BK006945.2| 613811 - INS T
 tpg|BK006949.2| 861091 + tpg|BK006949.2| 861210 - INS 
 tpg|BK006945.2| 525687 + tpg|BK006945.2| 525224 - INS 
 tpg|BK006945.2| 584248 + tpg|BK006945.2| 584106 - INS 
 tpg|BK006945.2| 53452 + tpg|BK006945.2| 53372 - INS 
 tpg|BK006949.2| 267710 + tpg|BK006949.2| 268435 - INS 
 tpg|BK006945.2| 1037926 + tpg|BK006945.2| 1037666 - INS 
 tpg|BK006945.2| 947271 + tpg|BK006945.2| 947013 - INS 
 tpg|BK006945.2| 727938 + tpg|BK006945.2| 727656 - INS 
 tpg|BK006949.2| 458225 + tpg|BK006949.2| 458709 - INS 
 tpg|BK006945.2| 401930 + tpg|BK006945.2| 401468 - INS 
 tpg|BK006945.2| 248694 + tpg|BK006945.2| 248718 - INS 
 tpg|BK006945.2| 581848 + tpg|BK006945.2| 581964 - INS 
 tpg|BK006945.2| 778568 + tpg|BK006945.2| 778691 - INS 
 tpg|BK006945.2| 393500 + tpg|BK006945.2| 393579 - INS 
 tpg|BK006945.2| 739197 + tpg|BK006945.2| 738772 - INS 
 tpg|BK006944.2| 650749 + tpg|BK006944.2| 651447 - INS 
 tpg|BK006945.2| 871967 + tpg|BK006945.2| 871481 - INS 
 tpg|BK006945.2| 1037245 + tpg|BK006945.2| 1036877 - INS 
 tpg|BK006945.2| 896705 + tpg|BK006945.2| 896889 - INS 
 tpg|BK006945.2| 583823 + tpg|BK006945.2| 583462 - INS 
 tpg|BK006945.2| 339038 + tpg|BK006945.2| 338495 - INS 
 tpg|BK006945.2| 851871 + tpg|BK006945.2| 851822 - INS 
 tpg|BK006945.2| 708688 + tpg|BK006945.2| 708296 - INS 
 tpg|BK006945.2| 56054 + tpg|BK006945.2| 55687 - INS 
 tpg|BK006945.2| 845518 + tpg|BK006945.2| tpg|BK006944.2| 845846 - INS 
 tpg|BK006945.2| 845518 + tpg|BK006945.2| tpg|BK006944.2| 845846 - INS 
638936 + tpg|BK006944.2| 639035 - INS 
 tpg|BK006945.2| 1005847 + tpg|BK006945.2| 1005612 - INS 
 tpg|BK006945.2| 510169 + tpg|BK006945.2| 510646 - INS 
 tpg|BK006944.2| 636673 + tpg|BK006944.2| 636681 - INS 
 tpg|BK006944.2| 77784 + tpg|BK006944.2| 77487 - INS 
 tpg|BK006949.2| 742892 + tpg|BK006949.2| 742601 - INS 
 tpg|BK006944.2| 280197 + tpg|BK006944.2| 280088 - INS 
 tpg|BK006949.2| 426685 + tpg|BK006949.2| 426061 - INS 
 tpg|BK006944.2| 279420 + tpg|BK006944.2| 279113 - INS 
 tpg|BK006944.2| 241491 + tpg|BK006944.2| 241546 - INS 
 tpg|BK006945.2| 375670 + tpg|BK006945.2| 375774 - INS 
 tpg|BK006944.2| 61335 + tpg|BK006944.2| 61546 - INS 
 tpg|BK006949.2| 110726 + tpg|BK006949.2| 110436 - INS 
 tpg|BK006945.2| 515024 + tpg|BK006945.2| 514860 - INS 
 tpg|BK006945.2| 37380 + tpg|BK006945.2| 37554 - INS 
 tpg|BK006944.2| 423127 + tpg|BK006944.2| 422613 - INS 
 tpg|BK006949.2| 504141 + tpg|BK006949.2| 503379 - INS 
 tpg|BK006945.2| 636375 + tpg|BK006945.2| 635670 - INS 
 tpg|BK006945.2| 749876 + tpg|BK006945.2| 750092 - INS 
 tpg|BK006945.2| 207139 + tpg|BK006945.2| 206895 - INS 
 tpg|BK006949.2| 919667 + tpg|BK006949.2| 919798 - INS GA
 tpg|BK006945.2| 889359 + tpg|BK006945.2| 888868 - INS 
 tpg|BK006945.2| 948860 + tpg|BK006945.2| 948510 - INS 
 tpg|BK006945.2| 332127 + tpg|BK006945.2| 332510 - INS 
 tpg|BK006945.2| 951504 + tpg|BK006945.2| 951927 - INS 
 tpg|BK006949.2| 718667 + tpg|BK006949.2| 717899 - INS 
 tpg|BK006945.2| 188100 + tpg|BK006945.2| 187802 - INS 
 tpg|BK006944.2| 493299 + tpg|BK006944.2| 492873 - INS 
 tpg|BK006945.2| 616107 + tpg|BK006945.2| 616807 - INS 
 tpg|BK006945.2| 414165 + tpg|BK006945.2| 413981 - INS 
 tpg|BK006945.2| 936964 + tpg|BK006945.2| 937413 - INS 
 tpg|BK006949.2| 756018 + tpg|BK006949.2| 755943 - INS 
 tpg|BK006945.2| 556235 + tpg|BK006945.2| 556257 - INS 
 tpg|BK006944.2| 505343 + tpg|BK006944.2| 505709 - INS TTATAACTTACAT
 tpg|BK006949.2| 659742 + tpg|BK006949.2| 660037 - INS 
 tpg|BK006945.2| 247238 + tpg|BK006945.2| 246519 - INS 
 tpg|BK006945.2| 806637 + tpg|BK006945.2| 806360 - INS 
 tpg|BK006944.2| 510666 + tpg|BK006944.2| 511382 - INS 
 tpg|BK006945.2| 133868 + tpg|BK006945.2| 133666 - INS 
 tpg|BK006945.2| 766810 + tpg|BK006945.2| 766856 - INS 
 tpg|BK006944.2| 297848 + tpg|BK006944.2| 297361 - INS 
 tpg|BK006945.2| 401308 + tpg|BK006945.2| 400625 - INS 
 tpg|BK006945.2| 615688 + tpg|BK006945.2| 615742 - INS 
 tpg|BK006945.2| 128346 + tpg|BK006945.2| 128496 - INS 
 tpg|BK006944.2| 82763 + tpg|BK006944.2| 82349 - INS 
 tpg|BK006945.2| 185764 + tpg|BK006945.2| 186105 - INS 
 tpg|BK006945.2| 516031 + tpg|BK006945.2| 515641 - INS 
 tpg|BK006945.2| 672985 + tpg|BK006945.2| 673061 - INS 
 tpg|BK006944.2| 558938 + tpg|BK006944.2| 559664 - INS 
 tpg|BK006945.2| 93887 + tpg|BK006945.2| 93460 - INS 
 tpg|BK006945.2| 22415 + tpg|BK006945.2| 22550 - INS 
 tpg|BK006945.2| 563914 + tpg|BK006945.2| 563716 - INS 
 tpg|BK006945.2| 667215 + tpg|BK006945.2| 666918 - INS 
 tpg|BK006945.2| 1022247 + tpg|BK006945.2| 1022118 - INS 
 tpg|BK006944.2| 657257 + tpg|BK006944.2| 657163 - INS 
 tpg|BK006945.2| 1051514 + tpg|BK006945.2| 1051130 - INS 
 tpg|BK006945.2| 361497 + tpg|BK006945.2| 361491 - INS 
 tpg|BK006945.2| 714142 + tpg|BK006945.2| 714341 - INS 
 tpg|BK006945.2| 929687 + tpg|BK006945.2| 929632 - INS 
 tpg|BK006945.2| 75778 + tpg|BK006945.2| 75444 - INS 
 tpg|BK006945.2| 651241 + tpg|BK006945.2| 651012 - INS 
 tpg|BK006945.2| 780650 + tpg|BK006945.2| 780551 - INS 
 tpg|BK006945.2| 135659 + tpg|BK006945.2| 136041 - INS 
 tpg|BK006945.2| 445905 + tpg|BK006945.2| 445830 - INS 
 tpg|BK006945.2| 831554 + tpg|BK006945.2| 831520 - INS 
 tpg|BK006945.2| 264850 + tpg|BK006945.2| 264966 - INS 
 tpg|BK006945.2| 342928 + tpg|BK006945.2| 342242 - INS 
 tpg|BK006944.2| 25651 + tpg|BK006944.2| 25734 - INS 
 tpg|BK006949.2| 705120 + tpg|BK006949.2| 705154 - INS 
 tpg|BK006949.2| 131618 + tpg|BK006949.2| 131581 - INS 
 tpg|BK006944.2| 177141 + tpg|BK006944.2| 176445 - INS 
 tpg|BK006949.2| 98784 + tpg|BK006949.2| 98575 - INS 
 tpg|BK006944.2| 178088 + tpg|BK006944.2| 177341 - INS 
 tpg|BK006944.2| 632361 + tpg|BK006944.2| 631591 - INS 
 tpg|BK006949.2| 46452 + tpg|BK006949.2| 46630 - INS 
 tpg|BK006944.2| 138660 + tpg|BK006944.2| 139249 - INS 
 tpg|BK006944.2| 130449 + tpg|BK006944.2| 130617 - INS 
 tpg|BK006949.2| 535184 + tpg|BK006949.2| 535169 - INS 
 tpg|BK006944.2| 106512 + tpg|BK006944.2| 105792 - INS 
 tpg|BK006949.2| 483922 + tpg|BK006949.2| 483184 - INS 
 tpg|BK006944.2| 514423 + tpg|BK006944.2| 514145 - INS 
 tpg|BK006944.2| 370549 + tpg|BK006944.2| 370709 - INS 
 tpg|BK006949.2| 565933 + tpg|BK006949.2| 565315 - INS 
 tpg|BK006944.2| 191229 + tpg|BK006944.2| 191025 - INS 
 tpg|BK006949.2| 256656 + tpg|BK006949.2| 257063 - INS 
 tpg|BK006944.2| 330934 + tpg|BK006944.2| 330718 - INS 
 tpg|BK006944.2| 544750 + tpg|BK006944.2| 544104 - INS 
 tpg|BK006944.2| 102027 + tpg|BK006944.2| 102730 - INS 
 tpg|BK006949.2| 101054 + tpg|BK006949.2| 100284 - INS 
 tpg|BK006944.2| 209601 + tpg|BK006944.2| 209033 - INS 
 tpg|BK006949.2| 530354 + tpg|BK006949.2| 530368 - INS 
 tpg|BK006949.2| 176830 + tpg|BK006949.2| 177227 - INS 
 tpg|BK006949.2| 903528 + tpg|BK006949.2| 903716 - INS 
 tpg|BK006949.2| 446563 + tpg|BK006949.2| 445868 - INS 
 tpg|BK006944.2| 201650 + tpg|BK006944.2| 202150 - INS 
 tpg|BK006949.2| 836610 + tpg|BK006949.2| 836134 - INS 
 tpg|BK006949.2| 550454 + tpg|BK006949.2| 549860 - INS 
 tpg|BK006944.2| 606293 + tpg|BK006944.2| 605715 - INS 
 tpg|BK006949.2| 636739 + tpg|BK006949.2| 637337 - INS 
 tpg|BK006949.2| 801951 + tpg|BK006949.2| 802590 - INS 
 tpg|BK006949.2| 244283 + tpg|BK006949.2| 244101 - INS 
 tpg|BK006944.2| 584259 + tpg|BK006944.2| 584109 - INS 
 tpg|BK006944.2| 599147 + tpg|BK006944.2| 599271 - INS 
 tpg|BK006949.2| 817342 + tpg|BK006949.2| 816959 - INS 
 tpg|BK006944.2| 641051 + tpg|BK006944.2| 640792 - INS 
 tpg|BK006944.2| 489774 + tpg|BK006944.2| 490078 - INS 
 tpg|BK006944.2| 212946 + tpg|BK006944.2| 212447 - INS 
 tpg|BK006949.2| 137138 + tpg|BK006949.2| 137686 - INS 
 tpg|BK006944.2| 648531 + tpg|BK006944.2| 648976 - INS 
 tpg|BK006944.2| 207215 + tpg|BK006944.2| 207328 - INS 
 tpg|BK006949.2| 308938 + tpg|BK006949.2| 309100 - INS 
 tpg|BK006944.2| 336016 + tpg|BK006944.2| 336180 - INS 
 tpg|BK006949.2| 735379 + tpg|BK006949.2| 734893 - INS 
 tpg|BK006949.2| 282923 + tpg|BK006949.2| 282552 - INS 
 tpg|BK006949.2| 796916 + tpg|BK006949.2| 796163 - INS 
 tpg|BK006944.2| 200965 + tpg|BK006944.2| 201256 - INS 
 tpg|BK006944.2| 51715 + tpg|BK006944.2| 51218 - INS 
 tpg|BK006949.2| 41638 + tpg|BK006949.2| 41604 - INS 
 tpg|BK006949.2| 113584 + tpg|BK006949.2| 113738 - INS 
 tpg|BK006944.2| 218787 + tpg|BK006944.2| 218819 - INS 
 tpg|BK006949.2| 905471 + tpg|BK006949.2| 905007 - INS 
 tpg|BK006949.2| 580663 + tpg|BK006949.2| 579938 - INS 
 tpg|BK006944.2| 72023 + tpg|BK006944.2| 72578 - INS 
 tpg|BK006944.2| 615879 + tpg|BK006944.2| 615404 - INS 
 tpg|BK006949.2| 620101 + tpg|BK006949.2| 620359 - INS 
 tpg|BK006944.2| 264322 + tpg|BK006944.2| 264170 - INS 
 tpg|BK006949.2| 681783 + tpg|BK006949.2| 681246 - INS 
 tpg|BK006944.2| 553151 + tpg|BK006944.2| 552754 - INS 
 tpg|BK006949.2| 712884 + tpg|BK006949.2| 712443 - INS 
 tpg|BK006944.2| 125396 + tpg|BK006944.2| 126133 - INS 
 tpg|BK006949.2| 302399 + tpg|BK006949.2| 302434 - INS 
 tpg|BK006944.2| 79005 + tpg|BK006944.2| 79204 - INS 
 tpg|BK006949.2| 526987 + tpg|BK006949.2| 526651 - INS 
 tpg|BK006944.2| 165975 + tpg|BK006944.2| 165572 - INS 
 tpg|BK006949.2| 172630 + tpg|BK006949.2| 172161 - INS 
 tpg|BK006944.2| 29591 + tpg|BK006944.2| 30154 - INS 
 tpg|BK006949.2| 104218 + tpg|BK006949.2| 104733 - INS 
 tpg|BK006944.2| 148365 + tpg|BK006944.2| 148027 - INS 
 tpg|BK006949.2| 478272 + tpg|BK006949.2| 477739 - INS 
 tpg|BK006944.2| 395354 + tpg|BK006944.2| 395053 - INS 
 tpg|BK006949.2| 102457 + tpg|BK006949.2| 102133 - INS 
 tpg|BK006944.2| 438367 + tpg|BK006944.2| 437612 - INS 
 tpg|BK006949.2| 162346 + tpg|BK006949.2| 161782 - INS 
 tpg|BK006944.2| 591167 + tpg|BK006944.2| 590707 - INS 
 tpg|BK006944.2| 590415 + tpg|BK006944.2| 590218 - INS 
 tpg|BK006944.2| 315937 + tpg|BK006944.2| 315967 - INS 
 tpg|BK006949.2| 900657 + tpg|BK006949.2| 900605 - INS 
 tpg|BK006944.2| 596133 + tpg|BK006944.2| 596841 - INS 
 tpg|BK006949.2| 127834 + tpg|BK006949.2| 128577 - INS 
 tpg|BK006944.2| 4957 + tpg|BK006944.2| 5416 - INS 
 tpg|BK006944.2| 112736 + tpg|BK006944.2| 112843 - INS 
 tpg|BK006949.2| 391389 + tpg|BK006949.2| 391097 - INS 
 tpg|BK006949.2| 367892 + tpg|BK006949.2| 367476 - INS 
 tpg|BK006949.2| 369498 + tpg|BK006949.2| 369645 - INS 
 tpg|BK006949.2| 249124 + tpg|BK006949.2| 248584 - INS 
 tpg|BK006944.2| 665487 + tpg|BK006944.2| 666220 - INS 
 tpg|BK006949.2| 614043 + tpg|BK006949.2| 614429 - INS 
 tpg|BK006944.2| 604063 + tpg|BK006944.2| 603400 - INS 
 tpg|BK006949.2| 784462 + tpg|BK006949.2| 784432 - INS 
 tpg|BK006944.2| 501978 + tpg|BK006944.2| 502739 - INS 
 tpg|BK006949.2| 389020 + tpg|BK006949.2| 388254 - INS 
 tpg|BK006944.2| 433842 + tpg|BK006944.2| 434013 - INS 
 tpg|BK006949.2| 47805 + tpg|BK006949.2| 47569 - INS 
 tpg|BK006949.2| 84933 + tpg|BK006949.2| 84863 - INS 
 tpg|BK006944.2| 509840 + tpg|BK006944.2| 509635 - INS 
 tpg|BK006949.2| 294321 + tpg|BK006949.2| 294557 - INS 
 tpg|BK006944.2| 103839 + tpg|BK006944.2| 103521 - INS 
 tpg|BK006949.2| 306341 + tpg|BK006949.2| 306265 - INS 
 tpg|BK006949.2| 295752 + tpg|BK006949.2| 295647 - INS 
 tpg|BK006944.2| 268780 + tpg|BK006944.2| 268646 - INS 
 tpg|BK006949.2| 463067 + tpg|BK006949.2| 462764 - INS 
 tpg|BK006944.2| 33925 + tpg|BK006944.2| 33195 - INS 
 tpg|BK006944.2| 634540 + tpg|BK006944.2| 635081 - INS 
 tpg|BK006949.2| 476130 + tpg|BK006949.2| 476036 - INS 
 tpg|BK006944.2| 565336 + tpg|BK006944.2| 565213 - INS 
 tpg|BK006944.2| 277971 + tpg|BK006944.2| 277528 - INS 
 tpg|BK006949.2| 583324 + tpg|BK006949.2| 583011 - INS 
 tpg|BK006944.2| 352197 + tpg|BK006944.2| 352037 - INS 
 tpg|BK006944.2| 233197 + tpg|BK006944.2| 233553 - INS 
 tpg|BK006949.2| 656440 + tpg|BK006949.2| 656582 - INS 
 tpg|BK006944.2| 403345 + tpg|BK006944.2| 403275 - INS 
 tpg|BK006944.2| 654402 + tpg|BK006944.2| 654103 - INS 
 tpg|BK006944.2| 390219 + tpg|BK006944.2| 389855 - INS 
 tpg|BK006944.2| 118133 + tpg|BK006944.2| 117740 - INS 
 tpg|BK006944.2| 113752 + tpg|BK006944.2| 113822 - INS 
 tpg|BK006949.2| 262687 + tpg|BK006949.2| 262939 - INS 
 tpg|BK006944.2| 491126 + tpg|BK006944.2| 491665 - INS 
 tpg|BK006944.2| 586982 + tpg|BK006944.2| 586985 - INS 
 tpg|BK006949.2| 666891 + tpg|BK006949.2| 666312 - INS 
 tpg|BK006944.2| 359097 + tpg|BK006944.2| 359306 - INS 
 tpg|BK006944.2| 320025 + tpg|BK006944.2| 319438 - INS 
 tpg|BK006949.2| 607866 + tpg|BK006949.2| 608585 - INS 
 tpg|BK006949.2| 911997 + tpg|BK006949.2| 911573 - INS 
 tpg|BK006944.2| 642165 + tpg|BK006944.2| 641936 - INS 
 tpg|BK006949.2| 115855 + tpg|BK006949.2| 115705 - INS 
 tpg|BK006944.2| 399936 + tpg|BK006944.2| 400481 - INS 
 tpg|BK006949.2| 141816 + tpg|BK006949.2| 141368 - INS 
 tpg|BK006944.2| 48919 + tpg|BK006944.2| 49414 - INS 
 tpg|BK006949.2| 556826 + tpg|BK006949.2| 556247 - INS 
 tpg|BK006944.2| 444079 + tpg|BK006944.2| 444012 - INS 
 tpg|BK006949.2| 189474 + tpg|BK006949.2| 188926 - INS 
 tpg|BK006949.2| 229943 + tpg|BK006949.2| 230594 - INS 
 tpg|BK006949.2| 669133 + tpg|BK006949.2| 669872 - INS 
 tpg|BK006944.2| 98453 + tpg|BK006944.2| 98469 - INS 
 tpg|BK006944.2| 289751 + tpg|BK006944.2| 289884 - INS 
 tpg|BK006949.2| 630826 + tpg|BK006949.2| 631354 - INS 
 tpg|BK006944.2| 84794 + tpg|BK006944.2| 84451 - INS 
 tpg|BK006949.2| 536808 + tpg|BK006949.2| 536492 - INS 
 tpg|BK006944.2| 228719 + tpg|BK006944.2| 228424 - INS 
 tpg|BK006944.2| 652527 + tpg|BK006944.2| 652750 - INS 
 tpg|BK006949.2| 926447 + tpg|BK006949.2| 926376 - INS 
 tpg|BK006944.2| 649961 + tpg|BK006944.2| 649635 - INS 
 tpg|BK006949.2| 720228 + tpg|BK006949.2| 719999 - INS 
 tpg|BK006944.2| 274345 + tpg|BK006944.2| 274314 - INS 
 tpg|BK006949.2| 485026 + tpg|BK006949.2| 485699 - INS 
 tpg|BK006944.2| 269873 + tpg|BK006944.2| 269573 - INS 
 tpg|BK006944.2| 567768 + tpg|BK006944.2| 568405 - INS 
 tpg|BK006949.2| 435423 + tpg|BK006949.2| 435445 - INS 
 tpg|BK006944.2| 71264 + tpg|BK006944.2| 70593 - INS 
 tpg|BK006949.2| 771554 + tpg|BK006949.2| 771588 - INS 
 tpg|BK006944.2| 65695 + tpg|BK006944.2| 65686 - INS 
 tpg|BK006949.2| 779215 + tpg|BK006949.2| 778988 - INS 
 tpg|BK006944.2| 231488 + tpg|BK006944.2| 230944 - INS 
 tpg|BK006949.2| 428222 + tpg|BK006949.2| 428188 - INS 
 tpg|BK006944.2| 609564 + tpg|BK006944.2| 610333 - INS 
 tpg|BK006949.2| 427414 + tpg|BK006949.2| 426912 - INS 
 tpg|BK006944.2| 387164 + tpg|BK006944.2| 387590 - INS 
 tpg|BK006949.2| 126045 + tpg|BK006949.2| 125567 - INS 
 tpg|BK006944.2| 433159 + tpg|BK006944.2| 432684 - INS 
 tpg|BK006949.2| 207561 + tpg|BK006949.2| 207428 - INS 
 tpg|BK006949.2| 581338 + tpg|BK006949.2| 580729 - INS 
 tpg|BK006944.2| 312223 + tpg|BK006944.2| 312773 - INS 
 tpg|BK006949.2| 602700 + tpg|BK006949.2| 603070 - INS 
 tpg|BK006944.2| 99985 + tpg|BK006944.2| 99867 - INS 
 tpg|BK006949.2| 276529 + tpg|BK006949.2| 276768 - INS 
 tpg|BK006944.2| 166998 + tpg|BK006944.2| 167756 - INS 
 tpg|BK006944.2| 235181 + tpg|BK006944.2| 234791 - INS 
 tpg|BK006949.2| 693834 + tpg|BK006949.2| 693074 - INS 
 tpg|BK006944.2| 233652 + tpg|BK006944.2| 234082 - INS 
 tpg|BK006949.2| 86066 + tpg|BK006949.2| 86579 - INS 
 tpg|BK006944.2| 431346 + tpg|BK006944.2| 431794 - INS 
 tpg|BK006949.2| 617829 + tpg|BK006949.2| 617268 - INS 
 tpg|BK006944.2| 157489 + tpg|BK006944.2| 156793 - INS 
 tpg|BK006944.2| 626091 + tpg|BK006944.2| 626013 - INS 
 tpg|BK006949.2| 222361 + tpg|BK006949.2| 221688 - INS 
 tpg|BK006949.2| 65918 + tpg|BK006949.2| 65534 - INS 
 tpg|BK006949.2| 585334 + tpg|BK006949.2| 584736 - INS 
 tpg|BK006944.2| 186689 + tpg|BK006944.2| 186866 - INS 
 tpg|BK006949.2| 932679 + tpg|BK006949.2| 932002 - INS 
 tpg|BK006944.2| 46982 + tpg|BK006944.2| 46439 - INS 
 tpg|BK006949.2| 20779 + tpg|BK006949.2| 20339 - INS 
 tpg|BK006949.2| 740419 + tpg|BK006949.2| 741029 - INS 
 tpg|BK006944.2| 545884 + tpg|BK006944.2| 545901 - INS 
 tpg|BK006944.2| 85756 + tpg|BK006944.2| 86435 - INS 
 tpg|BK006949.2| 291480 + tpg|BK006949.2| 291268 - INS 
 tpg|BK006944.2| 285319 + tpg|BK006944.2| 285354 - INS 
 tpg|BK006944.2| 90748 + tpg|BK006944.2| 90458 - INS 
 tpg|BK006949.2| 288715 + tpg|BK006949.2| 288386 - INS 
 tpg|BK006944.2| 523284 + tpg|BK006944.2| 522919 - INS 
 tpg|BK006949.2| 40782 + tpg|BK006949.2| 40166 - INS 
 tpg|BK006949.2| 124733 + tpg|BK006949.2| 124222 - INS 
 tpg|BK006949.2| 646404 + tpg|BK006949.2| 646553 - INS 
 tpg|BK006949.2| 27484 + tpg|BK006949.2| 27299 - INS 
 tpg|BK006949.2| 208994 + tpg|BK006949.2| 209245 - INS 
 tpg|BK006949.2| 795046 + tpg|BK006949.2| 794514 - INS 
 tpg|BK006949.2| 644672 + tpg|BK006949.2| 644097 - INS 
 tpg|BK006944.2| 127317 + tpg|BK006944.2| 127253 - INS 
 tpg|BK006949.2| 517426 + tpg|BK006949.2| 516979 - INS 
 tpg|BK006944.2| 253340 + tpg|BK006944.2| 252680 - INS 
 tpg|BK006944.2| 195822 + tpg|BK006944.2| 195482 - INS 
 tpg|BK006949.2| 672896 + tpg|BK006949.2| 672234 - INS 
 tpg|BK006944.2| 421306 + tpg|BK006944.2| 420865 - INS 
 tpg|BK006949.2| 335132 + tpg|BK006949.2| 334456 - INS 
 tpg|BK006944.2| 371943 + tpg|BK006944.2| 371498 - INS 
 tpg|BK006949.2| 432655 + tpg|BK006949.2| 432054 - INS 
 tpg|BK006944.2| 449915 + tpg|BK006944.2| 449578 - INS 
 tpg|BK006949.2| 240030 + tpg|BK006949.2| 239394 - INS 
 tpg|BK006944.2| 172070 + tpg|BK006944.2| 171668 - INS 
 tpg|BK006949.2| 563082 + tpg|BK006949.2| 562947 - INS 
 tpg|BK006944.2| 74717 + tpg|BK006944.2| 73982 - INS 
 tpg|BK006944.2| 368008 + tpg|BK006944.2| 367923 - INS 
 tpg|BK006949.2| 554060 + tpg|BK006949.2| 553646 - INS 
 tpg|BK006944.2| 287764 + tpg|BK006944.2| 287468 - INS 
 tpg|BK006949.2| 541600 + tpg|BK006949.2| 541500 - INS 
 tpg|BK006944.2| 577144 + tpg|BK006944.2| 577513 - INS 
 tpg|BK006944.2| 184572 + tpg|BK006944.2| 184330 - INS 
 tpg|BK006944.2| 13281 + tpg|BK006944.2| 13082 - INS 
 tpg|BK006949.2| 533220 + tpg|BK006949.2| 533825 - INS 
 tpg|BK006944.2| 323638 + tpg|BK006944.2| 324015 - INS 
 tpg|BK006949.2| 54107 + tpg|BK006949.2| 54786 - INS 
 tpg|BK006949.2| 460182 + tpg|BK006949.2| 459975 - INS 
 tpg|BK006949.2| 453941 + tpg|BK006949.2| 454013 - INS 
 tpg|BK006944.2| 216375 + tpg|BK006944.2| 216090 - INS 
 tpg|BK006949.2| 736160 + tpg|BK006949.2| 735742 - INS 
 tpg|BK006944.2| 83553 + tpg|BK006944.2| 83757 - INS 
 tpg|BK006949.2| 626169 + tpg|BK006949.2| 626342 - INS 
 tpg|BK006944.2| 575180 + tpg|BK006944.2| 575760 - INS 
 tpg|BK006944.2| 564436 + tpg|BK006944.2| 564271 - INS 
 tpg|BK006949.2| 404784 + tpg|BK006949.2| 405503 - INS 
 tpg|BK006944.2| 658341 + tpg|BK006944.2| 657922 - INS 
 tpg|BK006949.2| 235236 + tpg|BK006949.2| 234627 - INS 
 tpg|BK006944.2| 499862 + tpg|BK006944.2| 499122 - INS 
 tpg|BK006949.2| 233474 + tpg|BK006949.2| 233864 - INS 
 tpg|BK006949.2| 888432 + tpg|BK006949.2| 887878 - INS 
 tpg|BK006944.2| 137673 + tpg|BK006944.2| 136919 - INS 
 tpg|BK006949.2| 385188 + tpg|BK006949.2| 384479 - INS 
 tpg|BK006944.2| 227635 + tpg|BK006944.2| 226881 - INS 
 tpg|BK006944.2| 426152 + tpg|BK006944.2| 426747 - INS 
 tpg|BK006949.2| 887442 + tpg|BK006949.2| 887064 - INS 
 tpg|BK006944.2| 539341 + tpg|BK006944.2| 538661 - INS 
 tpg|BK006949.2| 103822 + tpg|BK006949.2| 103279 - INS 
 tpg|BK006944.2| 300778 + tpg|BK006944.2| 300335 - INS 
 tpg|BK006944.2| 32928 + tpg|BK006944.2| 32258 - INS 
 tpg|BK006949.2| 363449 + tpg|BK006949.2| 364115 - INS 
 tpg|BK006949.2| 599329 + tpg|BK006949.2| 598763 - INS 
 tpg|BK006944.2| 401975 + tpg|BK006944.2| 402168 - INS 
 tpg|BK006944.2| 150239 + tpg|BK006944.2| 149833 - INS 
 tpg|BK006949.2| 421533 + tpg|BK006949.2| 421205 - INS 
 tpg|BK006949.2| 612211 + tpg|BK006949.2| 612881 - INS 
 tpg|BK006944.2| 392881 + tpg|BK006944.2| 392905 - INS 
 tpg|BK006944.2| 613982 + tpg|BK006944.2| 613341 - INS 
 tpg|BK006949.2| 217058 + tpg|BK006949.2| 217559 - INS 
 tpg|BK006944.2| 145032 + tpg|BK006944.2| 144423 - INS 
 tpg|BK006944.2| 578557 + tpg|BK006944.2| 579151 - INS 
 tpg|BK006949.2| 520974 + tpg|BK006949.2| 520638 - INS 
 tpg|BK006944.2| 442250 + tpg|BK006944.2| 441745 - INS 
 tpg|BK006949.2| 592473 + tpg|BK006949.2| 592784 - INS 
 tpg|BK006949.2| 590147 + tpg|BK006949.2| 590589 - INS 
 tpg|BK006949.2| 239037 + tpg|BK006949.2| 238464 - INS 
 tpg|BK006949.2| 542404 + tpg|BK006949.2| 542585 - INS 
 tpg|BK006944.2| 484272 + tpg|BK006944.2| 484400 - INS 
 tpg|BK006949.2| 688114 + tpg|BK006949.2| 687844 - INS 
 tpg|BK006944.2| 627063 + tpg|BK006944.2| 626625 - INS 
 tpg|BK006949.2| 489462 + tpg|BK006949.2| 489525 - INS 
 tpg|BK006944.2| 24866 + tpg|BK006944.2| 24098 - INS 
 tpg|BK006949.2| 702792 + tpg|BK006949.2| 703336 - INS 
 tpg|BK006949.2| 89298 + tpg|BK006949.2| 88880 - INS 
 tpg|BK006944.2| 141562 + tpg|BK006944.2| 140939 - INS 
 tpg|BK006949.2| 134118 + tpg|BK006949.2| 134368 - INS 
 tpg|BK006944.2| 455514 + tpg|BK006944.2| 454845 - INS 
 tpg|BK006944.2| 353024 + tpg|BK006944.2| 352639 - INS 
 tpg|BK006944.2| 180662 + tpg|BK006944.2| 180738 - INS 
 tpg|BK006949.2| 772427 + tpg|BK006949.2| 772800 - INS 
 tpg|BK006944.2| 460202 + tpg|BK006944.2| 460026 - INS 
 tpg|BK006944.2| 502947 + tpg|BK006944.2| 503523 - INS T
 tpg|BK006944.2| 532902 + tpg|BK006944.2| 533046 - INS 
 tpg|BK006949.2| 270813 + tpg|BK006949.2| 271496 - INS 
 tpg|BK006944.2| 550474 + tpg|BK006944.2| 550226 - INS 
 tpg|BK006944.2| 128659 + tpg|BK006944.2| 128882 - INS 
 tpg|BK006949.2| 214674 + tpg|BK006949.2| 214443 - INS 
 tpg|BK006944.2| 166363 + tpg|BK006944.2| 166126 - INS 
 tpg|BK006944.2| 483655 + tpg|BK006944.2| 483050 - INS 
 tpg|BK006949.2| 655303 + tpg|BK006949.2| 654531 - INS 
 tpg|BK006944.2| 471894 + tpg|BK006944.2| 471602 - INS 
 tpg|BK006949.2| 216335 + tpg|BK006949.2| 216152 - INS 
 tpg|BK006944.2| 512342 + tpg|BK006944.2| 512208 - INS 
 tpg|BK006944.2| 526112 + tpg|BK006944.2| 526484 - INS 
 tpg|BK006949.2| 798820 + tpg|BK006949.2| 799510 - INS 
 tpg|BK006944.2| 406245 + tpg|BK006944.2| 406748 - INS 
 tpg|BK006949.2| 106639 + tpg|BK006949.2| 106068 - INS 
 tpg|BK006944.2| 388932 + tpg|BK006944.2| 388733 - INS 
 tpg|BK006944.2| 581895 + tpg|BK006944.2| 582525 - INS 
 tpg|BK006944.2| 192472 + tpg|BK006944.2| 192832 - INS 
 tpg|BK006944.2| 591630 + tpg|BK006944.2| 592320 - INS 
 tpg|BK006944.2| 190743 + tpg|BK006944.2| 190219 - INS 
 tpg|BK006944.2| 595374 + tpg|BK006944.2| 595352 - INS 
 tpg|BK006949.2| 539682 + tpg|BK006949.2| 538964 - INS 
 tpg|BK006949.2| 670885 + tpg|BK006949.2| 671436 - INS 
 tpg|BK006944.2| 1059 + tpg|BK006944.2| 827 - INS 
 tpg|BK006949.2| 338199 + tpg|BK006949.2| 337544 - INS 
 tpg|BK006944.2| 45118 + tpg|BK006944.2| 44516 - INS 
 tpg|BK006949.2| 21291 + tpg|BK006949.2| 20867 - INS 
 tpg|BK006944.2| 348558 + tpg|BK006944.2| 347927 - INS 
 tpg|BK006949.2| 468109 + tpg|BK006949.2| 468837 - INS 
 tpg|BK006949.2| 168323 + tpg|BK006949.2| 168086 - INS 
 tpg|BK006944.2| 347127 + tpg|BK006944.2| 346368 - INS 
 tpg|BK006949.2| 164178 + tpg|BK006949.2| 163645 - INS 
 tpg|BK006949.2| 44249 + tpg|BK006949.2| 43530 - INS 
 tpg|BK006944.2| 36380 + tpg|BK006944.2| 35657 - INS 
 tpg|BK006944.2| 48062 + tpg|BK006944.2| 48653 - INS 
 tpg|BK006944.2| 306495 + tpg|BK006944.2| 306362 - INS 
 tpg|BK006949.2| 338793 + tpg|BK006949.2| 338615 - INS 
 tpg|BK006944.2| 304321 + tpg|BK006944.2| 304239 - INS 
 tpg|BK006944.2| 408738 + tpg|BK006944.2| 409276 - INS 
 tpg|BK006944.2| 151767 + tpg|BK006944.2| 151993 - INS 
 tpg|BK006949.2| 292886 + tpg|BK006949.2| 292737 - INS 
 tpg|BK006944.2| 138216 + tpg|BK006944.2| 137633 - INS 
 tpg|BK006949.2| 151057 + tpg|BK006949.2| 151465 - INS 
 tpg|BK006944.2| 445986 + tpg|BK006944.2| 445330 - INS 
 tpg|BK006944.2| 236421 + tpg|BK006944.2| 236542 - INS 
 tpg|BK006944.2| 515054 + tpg|BK006944.2| 515104 - INS 
 tpg|BK006944.2| 508746 + tpg|BK006944.2| 508947 - INS 
 tpg|BK006949.2| 340632 + tpg|BK006949.2| 340300 - INS 
 tpg|BK006944.2| 562964 + tpg|BK006944.2| 563269 - INS 
 tpg|BK006944.2| 574684 + tpg|BK006944.2| 574369 - INS 
 tpg|BK006949.2| 723586 + tpg|BK006949.2| 723268 - INS 
 tpg|BK006944.2| 10982 + tpg|BK006944.2| 10810 - INS 
 tpg|BK006949.2| 724995 + tpg|BK006949.2| 725201 - INS 
 tpg|BK006944.2| 495084 + tpg|BK006944.2| 495476 - INS 
 tpg|BK006949.2| 940032 + tpg|BK006949.2| 939841 - INS 
 tpg|BK006944.2| 549051 + tpg|BK006944.2| 548733 - INS 
 tpg|BK006949.2| 783340 + tpg|BK006949.2| 783441 - INS 
 tpg|BK006944.2| 583361 + tpg|BK006944.2| 583278 - INS 
 tpg|BK006949.2| 114521 + tpg|BK006949.2| 115189 - INS 
 tpg|BK006944.2| 411496 + tpg|BK006944.2| 410895 - INS 
 tpg|BK006944.2| 410205 + tpg|BK006944.2| 409772 - INS 
 tpg|BK006949.2| 484324 + tpg|BK006949.2| 484165 - INS 
 tpg|BK006949.2| 325822 + tpg|BK006949.2| 325115 - INS 
 tpg|BK006944.2| 428594 + tpg|BK006944.2| 428441 - INS 
 tpg|BK006944.2| 430476 + tpg|BK006944.2| 430418 - INS 
 tpg|BK006944.2| 173598 + tpg|BK006944.2| 172983 - INS 
 tpg|BK006949.2| 436808 + tpg|BK006949.2| 436219 - INS 
 tpg|BK006944.2| 189414 + tpg|BK006944.2| 188674 - INS 
 tpg|BK006944.2| 364468 + tpg|BK006944.2| 364479 - INS 
 tpg|BK006949.2| 405989 + tpg|BK006949.2| 406157 - INS 
 tpg|BK006944.2| 248735 + tpg|BK006944.2| 249332 - INS 
 tpg|BK006949.2| 331251 + tpg|BK006949.2| 331710 - INS 
 tpg|BK006944.2| 42225 + tpg|BK006944.2| 42490 - INS 
 tpg|BK006944.2| 101675 + tpg|BK006944.2| 102290 - INS 
 tpg|BK006944.2| 416104 + tpg|BK006944.2| 415520 - INS 
 tpg|BK006949.2| 505609 + tpg|BK006949.2| 505596 - INS 
 tpg|BK006949.2| 782360 + tpg|BK006949.2| 782801 - INS 
 tpg|BK006944.2| 566826 + tpg|BK006944.2| 566608 - INS 
 tpg|BK006944.2| 259319 + tpg|BK006944.2| 258608 - INS 
 tpg|BK006944.2| 419484 + tpg|BK006944.2| 418967 - INS 
 tpg|BK006944.2| 106921 + tpg|BK006944.2| 107668 - INS 
 tpg|BK006949.2| 78863 + tpg|BK006949.2| 78175 - INS 
 tpg|BK006944.2| 571694 + tpg|BK006944.2| 571777 - INS 
 tpg|BK006944.2| 602352 + tpg|BK006944.2| 601889 - INS 
 tpg|BK006949.2| 870849 + tpg|BK006949.2| 870794 - INS 
 tpg|BK006944.2| 378784 + tpg|BK006944.2| 378463 - INS 
 tpg|BK006944.2| 473061 + tpg|BK006944.2| 472754 - INS 
 tpg|BK006944.2| 156575 + tpg|BK006944.2| 156086 - INS 
 tpg|BK006944.2| 456377 + tpg|BK006944.2| 456163 - INS 
 tpg|BK006949.2| 653810 + tpg|BK006949.2| 653496 - INS 
 tpg|BK006944.2| 539669 + tpg|BK006944.2| 539435 - INS 
 tpg|BK006949.2| 265777 + tpg|BK006949.2| 265725 - INS 
 tpg|BK006944.2| 542398 + tpg|BK006944.2| 542165 - INS 
 tpg|BK006949.2| 642060 + tpg|BK006949.2| 642358 - INS 
 tpg|BK006944.2| 425670 + tpg|BK006944.2| 426060 - INS 
 tpg|BK006949.2| 639833 + tpg|BK006949.2| 639988 - INS 
 tpg|BK006949.2| 150221 + tpg|BK006949.2| 149494 - INS 
 tpg|BK006944.2| 20145 + tpg|BK006944.2| 19701 - INS 
 tpg|BK006949.2| 355095 + tpg|BK006949.2| 355057 - INS 
 tpg|BK006944.2| 15226 + tpg|BK006944.2| 14772 - INS 
 tpg|BK006949.2| 250462 + tpg|BK006949.2| 250572 - INS 
 tpg|BK006944.2| 261691 + tpg|BK006944.2| 261821 - INS 
 tpg|BK006944.2| 254621 + tpg|BK006944.2| 254721 - INS 
 tpg|BK006949.2| 433598 + tpg|BK006949.2| 433776 - INS 
 tpg|BK006944.2| 109658 + tpg|BK006944.2| 110229 - INS 
 tpg|BK006944.2| 253786 + tpg|BK006944.2| 253680 - INS 
 tpg|BK006949.2| 629877 + tpg|BK006949.2| 629169 - INS 
 tpg|BK006944.2| 258017 + tpg|BK006944.2| 257416 - INS 
 tpg|BK006949.2| 77603 + tpg|BK006949.2| 76993 - INS 
 tpg|BK006944.2| 466969 + tpg|BK006944.2| 466702 - INS 
 tpg|BK006944.2| 523989 + tpg|BK006944.2| 524336 - INS 
 tpg|BK006944.2| 537794 + tpg|BK006944.2| 537534 - INS 
 tpg|BK006944.2| 225804 + tpg|BK006944.2| 225489 - INS 
 tpg|BK006949.2| 832359 + tpg|BK006949.2| 832072 - INS 
 tpg|BK006949.2| 495627 + tpg|BK006949.2| 495570 - INS 
 tpg|BK006944.2| 407898 + tpg|BK006944.2| 407506 - INS 
 tpg|BK006949.2| 260437 + tpg|BK006949.2| 260241 - INS 
 tpg|BK006944.2| 7436 + tpg|BK006944.2| 7010 - INS 
 tpg|BK006949.2| 461454 + tpg|BK006949.2| 461352 - INS 
 tpg|BK006944.2| 324823 + tpg|BK006944.2| 325412 - INS 
 tpg|BK006944.2| 204954 + tpg|BK006944.2| 204891 - INS 
 tpg|BK006944.2| 605363 + tpg|BK006944.2| 604965 - INS 
 tpg|BK006949.2| 390052 + tpg|BK006949.2| 389372 - INS 
 tpg|BK006944.2| 347714 + tpg|BK006944.2| 347118 - INS 
 tpg|BK006944.2| 42888 + tpg|BK006944.2| 43449 - INS 
 tpg|BK006949.2| 513610 + tpg|BK006949.2| 514197 - INS 
 tpg|BK006944.2| 326810 + tpg|BK006944.2| 327089 - INS 
 tpg|BK006944.2| 66841 + tpg|BK006944.2| 66553 - INS 
 tpg|BK006949.2| 696947 + tpg|BK006949.2| 696517 - INS 
 tpg|BK006944.2| 349283 + tpg|BK006944.2| 349682 - INS 
 tpg|BK006944.2| 70796 + tpg|BK006944.2| 70099 - INS 
 tpg|BK006944.2| 617473 + tpg|BK006944.2| 616963 - INS 
 tpg|BK006944.2| 344250 + tpg|BK006944.2| 343976 - INS 
 tpg|BK006949.2| 133531 + tpg|BK006949.2| 134017 - INS 
 tpg|BK006944.2| 295801 + tpg|BK006944.2| 295765 - INS 
 tpg|BK006949.2| 121683 + tpg|BK006949.2| 122134 - INS 
 tpg|BK006944.2| 62610 + tpg|BK006944.2| 62269 - INS 
 tpg|BK006944.2| 197846 + tpg|BK006944.2| 198438 - INS 
 tpg|BK006949.2| 142590 + tpg|BK006949.2| 142136 - INS 
 tpg|BK006944.2| 194504 + tpg|BK006944.2| 194076 - INS 
 tpg|BK006944.2| 413604 + tpg|BK006944.2| 413269 - INS 
 tpg|BK006944.2| 160561 + tpg|BK006944.2| 160599 - INS 
 tpg|BK006949.2| 175152 + tpg|BK006949.2| 174636 - INS 
 tpg|BK006944.2| 75566 + tpg|BK006944.2| 75118 - INS 
 tpg|BK006949.2| 122757 + tpg|BK006949.2| 122580 - INS 
 tpg|BK006944.2| 80389 + tpg|BK006944.2| 79678 - INS 
 tpg|BK006949.2| 127338 + tpg|BK006949.2| 126880 - INS 
 tpg|BK006944.2| 298285 + tpg|BK006944.2| 298120 - INS 
 tpg|BK006944.2| 470480 + tpg|BK006944.2| 470353 - INS 
 tpg|BK006944.2| 438889 + tpg|BK006944.2| 438741 - INS 
 tpg|BK006944.2| 618417 + tpg|BK006944.2| 617712 - INS 
 tpg|BK006944.2| 396057 + tpg|BK006944.2| 396041 - INS 
 tpg|BK006944.2| 247983 + tpg|BK006944.2| 247849 - INS 
 tpg|BK006944.2| 321667 + tpg|BK006944.2| 321203 - INS 
 tpg|BK006949.2| 769448 + tpg|BK006949.2| 769964 - INS 
 tpg|BK006944.2| 250258 + tpg|BK006944.2| 250279 - INS 
 tpg|BK006949.2| 350454 + tpg|BK006949.2| 350055 - INS 
 tpg|BK006944.2| 439537 + tpg|BK006944.2| 439584 - INS 
 tpg|BK006949.2| 67787 + tpg|BK006949.2| 67556 - INS 
 tpg|BK006944.2| 320534 + tpg|BK006944.2| 320255 - INS 
 tpg|BK006949.2| 824397 + tpg|BK006949.2| 824983 - INS 
 tpg|BK006944.2| 468151 + tpg|BK006944.2| 467792 - INS 
 tpg|BK006944.2| 232517 + tpg|BK006944.2| 232397 - INS 
 tpg|BK006949.2| 873476 + tpg|BK006949.2| 872771 - INS 
 tpg|BK006944.2| 391450 + tpg|BK006944.2| 391458 - INS 
 tpg|BK006944.2| 135759 + tpg|BK006944.2| 135473 - INS 
 tpg|BK006944.2| 55730 + tpg|BK006944.2| 56025 - INS 
 tpg|BK006944.2| 39290 + tpg|BK006944.2| 39354 - INS 
 tpg|BK006949.2| 203872 + tpg|BK006949.2| 203907 - INS 
 tpg|BK006944.2| 374900 + tpg|BK006944.2| 374358 - INS 
 tpg|BK006944.2| 551483 + tpg|BK006944.2| 551695 - INS 
 tpg|BK006944.2| 133454 + tpg|BK006944.2| 133015 - INS 
 tpg|BK006949.2| 201383 + tpg|BK006949.2| 201847 - INS 
 tpg|BK006944.2| 560760 + tpg|BK006944.2| 560702 - INS 
 tpg|BK006944.2| 476491 + tpg|BK006944.2| 476995 - INS 
 tpg|BK006949.2| 651847 + tpg|BK006949.2| 651398 - INS 
 tpg|BK006944.2| 237349 + tpg|BK006944.2| 237244 - INS 
 tpg|BK006944.2| 307727 + tpg|BK006944.2| 307315 - INS 
 tpg|BK006944.2| 607328 + tpg|BK006944.2| 607857 - INS 
 tpg|BK006949.2| 882763 + tpg|BK006949.2| 882392 - INS 
 tpg|BK006944.2| 354882 + tpg|BK006944.2| 354651 - INS 
 tpg|BK006944.2| 553828 + tpg|BK006944.2| 553631 - INS 
 tpg|BK006944.2| 174263 + tpg|BK006944.2| 173492 - INS 
 tpg|BK006944.2| 397090 + tpg|BK006944.2| 396631 - INS 
 tpg|BK006949.2| 548604 + tpg|BK006949.2| 549235 - INS 
 tpg|BK006944.2| 263320 + tpg|BK006944.2| 262921 - INS 
 tpg|BK006944.2| 51012 + tpg|BK006944.2| 50728 - INS 
 tpg|BK006949.2| 259400 + tpg|BK006949.2| 258751 - INS 
 tpg|BK006944.2| 517277 + tpg|BK006944.2| 516987 - INS 
 tpg|BK006944.2| 536697 + tpg|BK006944.2| 536506 - INS 
 tpg|BK006949.2| 707563 + tpg|BK006949.2| 707548 - INS 
 tpg|BK006944.2| 573715 + tpg|BK006944.2| 573497 - INS 
 tpg|BK006944.2| 436004 + tpg|BK006944.2| 436315 - INS 
 tpg|BK006949.2| 196555 + tpg|BK006949.2| 195965 - INS 
 tpg|BK006944.2| 546828 + tpg|BK006944.2| 547112 - INS 
 tpg|BK006944.2| 343510 + tpg|BK006944.2| 343429 - INS 
 tpg|BK006949.2| 192774 + tpg|BK006949.2| 192524 - INS 
 tpg|BK006944.2| 469387 + tpg|BK006944.2| 469333 - INS 
 tpg|BK006944.2| 501074 + tpg|BK006944.2| 500376 - INS 
 tpg|BK006944.2| 199310 + tpg|BK006944.2| 199306 - INS 
 tpg|BK006949.2| 674661 + tpg|BK006949.2| 673970 - INS 
 tpg|BK006944.2| 112055 + tpg|BK006944.2| 111989 - INS 
 tpg|BK006949.2| 897709 + tpg|BK006949.2| 898031 - INS 
 tpg|BK006944.2| 588186 + tpg|BK006944.2| 587695 - INS 
 tpg|BK006949.2| 178884 + tpg|BK006949.2| 179400 - INS 
 tpg|BK006944.2| 556439 + tpg|BK006944.2| 556491 - INS 
 tpg|BK006949.2| 893082 + tpg|BK006949.2| 893697 - INS 
 tpg|BK006944.2| 593097 + tpg|BK006944.2| 592796 - INS 
 tpg|BK006949.2| 279846 + tpg|BK006949.2| 279768 - INS 
 tpg|BK006944.2| 429615 + tpg|BK006944.2| 429664 - INS 
 tpg|BK006944.2| 606779 + tpg|BK006944.2| 606240 - INS 
 tpg|BK006944.2| 182602 + tpg|BK006944.2| 182975 - INS 
 tpg|BK006944.2| 67398 + tpg|BK006944.2| 67206 - INS 
 tpg|BK006944.2| 7927 + tpg|BK006944.2| 8636 - INS 
 tpg|BK006944.2| 353800 + tpg|BK006944.2| 353588 - INS 
 tpg|BK006944.2| 462053 + tpg|BK006944.2| 461864 - INS 
 tpg|BK006944.2| 333128 + tpg|BK006944.2| 333581 - INS 
 tpg|BK006944.2| 381028 + tpg|BK006944.2| 380656 - INS 
 tpg|BK006944.2| 588930 + tpg|BK006944.2| 588520 - INS 
 tpg|BK006944.2| 581041 + tpg|BK006944.2| 580365 - INS 
 tpg|BK006944.2| 18219 + tpg|BK006944.2| 18172 - INS 
 tpg|BK006944.2| 111508 + tpg|BK006944.2| 110799 - INS 
 tpg|BK006944.2| 123445 + tpg|BK006944.2| 123373 - INS 
 tpg|BK006944.2| 213413 + tpg|BK006944.2| 212995 - INS 
 tpg|BK006944.2| 611219 + tpg|BK006944.2| 611967 - INS 
 tpg|BK006944.2| 496951 + tpg|BK006944.2| 497254 - INS 
 tpg|BK006944.2| 38668 + tpg|BK006944.2| 38438 - INS 
 tpg|BK006944.2| 158282 + tpg|BK006944.2| 158845 - INS 
 tpg|BK006944.2| 342767 + tpg|BK006944.2| 342568 - INS 
 tpg|BK006944.2| 1972 + tpg|BK006944.2| 2304 - INS 
 tpg|BK006944.2| 175155 + tpg|BK006944.2| 174897 - INS 
 tpg|BK006944.2| 446519 + tpg|BK006944.2| 446261 - INS 
 tpg|BK006944.2| 644355 + tpg|BK006944.2| 645013 - INS 
 tpg|BK006944.2| 381558 + tpg|BK006944.2| 381224 - INS 
 tpg|BK006944.2| 485243 + tpg|BK006944.2| 484997 - INS 
 tpg|BK006944.2| 242743 + tpg|BK006944.2| 242289 - INS 
 tpg|BK006944.2| 662041 + tpg|BK006944.2| 661366 - INS 
 tpg|BK006949.2| 691460 + tpg|BK006949.2| 690953 - INS 
 tpg|BK006949.2| 296501 + tpg|BK006949.2| 296544 - INS 
 tpg|BK006949.2| 716429 + tpg|BK006949.2| 717163 - INS 
 tpg|BK006949.2| 385969 + tpg|BK006949.2| 386688 - INS 
 tpg|BK006949.2| 764780 + tpg|BK006949.2| 764707 - INS 
 tpg|BK006949.2| 895386 + tpg|BK006949.2| 895248 - INS 
 tpg|BK006949.2| 638703 + tpg|BK006949.2| 638771 - INS 
 tpg|BK006949.2| 330595 + tpg|BK006949.2| 330786 - INS 
 tpg|BK006949.2| 934533 + tpg|BK006949.2| 935078 - INS 
 tpg|BK006949.2| 859369 + tpg|BK006949.2| 858800 - INS 
 tpg|BK006949.2| 166826 + tpg|BK006949.2| 166742 - INS 
 tpg|BK006949.2| 377180 + tpg|BK006949.2| 376898 - INS 
 tpg|BK006949.2| 868781 + tpg|BK006949.2| 868031 - INS 
 tpg|BK006949.2| 237364 + tpg|BK006949.2| 236631 - INS 
 tpg|BK006949.2| 381595 + tpg|BK006949.2| 381421 - INS 
 tpg|BK006949.2| 793404 + tpg|BK006949.2| 792794 - INS 
 tpg|BK006949.2| 726910 + tpg|BK006949.2| 727008 - INS 
 tpg|BK006949.2| 204817 + tpg|BK006949.2| 205464 - INS 
 tpg|BK006949.2| 922255 + tpg|BK006949.2| 922006 - INS 
 tpg|BK006949.2| 155327 + tpg|BK006949.2| 155527 - INS 
 tpg|BK006949.2| 165051 + tpg|BK006949.2| 164367 - INS 
 tpg|BK006949.2| 169136 + tpg|BK006949.2| 168704 - INS 
 tpg|BK006949.2| 423060 + tpg|BK006949.2| 423030 - INS 
 tpg|BK006949.2| 173190 + tpg|BK006949.2| 173569 - INS 
 tpg|BK006949.2| 572257 + tpg|BK006949.2| 572950 - INS 
 tpg|BK006949.2| 575021 + tpg|BK006949.2| 575714 - INS 
 tpg|BK006949.2| 653049 + tpg|BK006949.2| 652736 - INS 
 tpg|BK006949.2| 192117 + tpg|BK006949.2| 191953 - INS 
 tpg|BK006949.2| 616983 + tpg|BK006949.2| 616577 - INS 
 tpg|BK006949.2| 823934 + tpg|BK006949.2| 823409 - INS 
 tpg|BK006949.2| 916510 + tpg|BK006949.2| 916096 - INS 
 tpg|BK006949.2| 697650 + tpg|BK006949.2| 698075 - INS 
 tpg|BK006949.2| 232778 + tpg|BK006949.2| 232542 - INS 
 tpg|BK006949.2| 246093 + tpg|BK006949.2| 245829 - INS 
 tpg|BK006949.2| 258578 + tpg|BK006949.2| 257874 - INS 
 tpg|BK006949.2| 497005 + tpg|BK006949.2| 496697 - INS 
 tpg|BK006949.2| 152386 + tpg|BK006949.2| 152278 - INS 
 tpg|BK006949.2| 53181 + tpg|BK006949.2| 53792 - INS 
 tpg|BK006949.2| 336384 + tpg|BK006949.2| 335850 - INS 
 tpg|BK006949.2| 182762 + tpg|BK006949.2| 182319 - INS 
 tpg|BK006949.2| 348451 + tpg|BK006949.2| 348334 - INS 
 tpg|BK006949.2| 792034 + tpg|BK006949.2| 791886 - INS 
 tpg|BK006949.2| 866963 + tpg|BK006949.2| 867262 - INS 
 tpg|BK006949.2| 649898 + tpg|BK006949.2| 649256 - INS 
 tpg|BK006949.2| 788331 + tpg|BK006949.2| 788164 - INS 
 tpg|BK006949.2| 264160 + tpg|BK006949.2| 263949 - INS 
 tpg|BK006949.2| 378494 + tpg|BK006949.2| 378126 - INS 
 tpg|BK006949.2| 22073 + tpg|BK006949.2| 22594 - INS 
 tpg|BK006949.2| 743499 + tpg|BK006949.2| 744042 - INS 
 tpg|BK006949.2| 615458 + tpg|BK006949.2| 615253 - INS 
 tpg|BK006949.2| 95707 + tpg|BK006949.2| 95627 - INS 
 tpg|BK006949.2| 480141 + tpg|BK006949.2| 479520 - INS 
 tpg|BK006949.2| 706216 + tpg|BK006949.2| 706603 - INS 
 tpg|BK006949.2| 775732 + tpg|BK006949.2| 774960 - INS 
 tpg|BK006949.2| 764392 + tpg|BK006949.2| 763970 - INS 
 tpg|BK006949.2| 380373 + tpg|BK006949.2| 379624 - INS 
 tpg|BK006949.2| 333292 + tpg|BK006949.2| 333165 - INS 
 tpg|BK006949.2| 424794 + tpg|BK006949.2| 424685 - INS 
 tpg|BK006949.2| 180728 + tpg|BK006949.2| 180359 - INS 
 tpg|BK006949.2| 229282 + tpg|BK006949.2| 229204 - INS 
 tpg|BK006949.2| 719762 + tpg|BK006949.2| 719376 - INS 
 tpg|BK006949.2| 543232 + tpg|BK006949.2| 543204 - INS 
 tpg|BK006949.2| 91285 + tpg|BK006949.2| 90967 - INS 
 tpg|BK006949.2| 327726 + tpg|BK006949.2| 327443 - INS 
 tpg|BK006949.2| 679099 + tpg|BK006949.2| 679650 - INS 
 tpg|BK006949.2| 658049 + tpg|BK006949.2| 658750 - INS 
 tpg|BK006949.2| 190627 + tpg|BK006949.2| 190066 - INS 
 tpg|BK006949.2| 190996 + tpg|BK006949.2| 191298 - INS 
 tpg|BK006949.2| 314493 + tpg|BK006949.2| 314464 - INS 
 tpg|BK006949.2| 220731 + tpg|BK006949.2| 220451 - INS 
 tpg|BK006949.2| 299760 + tpg|BK006949.2| 299178 - INS 
 tpg|BK006949.2| 591719 + tpg|BK006949.2| 591345 - INS 
 tpg|BK006949.2| 570834 + tpg|BK006949.2| 570658 - INS 
 tpg|BK006949.2| 607431 + tpg|BK006949.2| 606956 - INS 
 tpg|BK006949.2| 246830 + tpg|BK006949.2| 246814 - INS 
 tpg|BK006949.2| 610199 + tpg|BK006949.2| 610128 - INS 
 tpg|BK006949.2| 482099 + tpg|BK006949.2| 482393 - INS 
 tpg|BK006949.2| 561291 + tpg|BK006949.2| 562033 - INS 
 tpg|BK006949.2| 281130 + tpg|BK006949.2| 280675 - INS 
 tpg|BK006949.2| 917667 + tpg|BK006949.2| 917076 - INS 
 tpg|BK006949.2| 49726 + tpg|BK006949.2| 49844 - INS 
 tpg|BK006949.2| 492519 + tpg|BK006949.2| 491805 - INS 
 tpg|BK006949.2| 551139 + tpg|BK006949.2| 551599 - INS 
 tpg|BK006949.2| 275877 + tpg|BK006949.2| 275626 - INS 
 tpg|BK006949.2| 912687 + tpg|BK006949.2| 912109 - INS 
 tpg|BK006949.2| 927595 + tpg|BK006949.2| 927047 - INS 
 tpg|BK006949.2| 694522 + tpg|BK006949.2| 694470 - INS 
 tpg|BK006949.2| 695841 + tpg|BK006949.2| 695468 - INS 
 tpg|BK006949.2| 710991 + tpg|BK006949.2| 710854 - INS 
 tpg|BK006949.2| 154359 + tpg|BK006949.2| 154321 - INS 
 tpg|BK006949.2| 298046 + tpg|BK006949.2| 297760 - INS 
 tpg|BK006949.2| 715757 + tpg|BK006949.2| 715793 - INS 
 tpg|BK006949.2| 148590 + tpg|BK006949.2| 148506 - INS 
 tpg|BK006949.2| 117509 + tpg|BK006949.2| 117490 - INS 
 tpg|BK006949.2| 875965 + tpg|BK006949.2| 876664 - INS 
 tpg|BK006949.2| 17839 + tpg|BK006949.2| 17145 - INS 
 tpg|BK006949.2| 394963 + tpg|BK006949.2| 394837 - INS 
 tpg|BK006949.2| 869952 + tpg|BK006949.2| 870403 - INS 
 tpg|BK006949.2| 359561 + tpg|BK006949.2| 359942 - INS 
 tpg|BK006949.2| 843469 + tpg|BK006949.2| 842839 - INS 
 tpg|BK006949.2| 371528 + tpg|BK006949.2| 370934 - INS 
 tpg|BK006949.2| 134548 + tpg|BK006949.2| 135321 - INS 
 tpg|BK006949.2| 746222 + tpg|BK006949.2| 745904 - INS 
 tpg|BK006949.2| 143003 + tpg|BK006949.2| 142836 - INS 
 tpg|BK006949.2| 32621 + tpg|BK006949.2| 32274 - INS 
 tpg|BK006949.2| 597098 + tpg|BK006949.2| 597527 - INS 
 tpg|BK006949.2| 107549 + tpg|BK006949.2| 106850 - INS 
 tpg|BK006949.2| 554843 + tpg|BK006949.2| 554318 - INS 
 tpg|BK006949.2| 713401 + tpg|BK006949.2| 713332 - INS 
 tpg|BK006949.2| 772926 + tpg|BK006949.2| 773616 - INS 
 tpg|BK006949.2| 352470 + tpg|BK006949.2| 353042 - INS 
 tpg|BK006949.2| 766196 + tpg|BK006949.2| 765584 - INS 
 tpg|BK006949.2| 449248 + tpg|BK006949.2| 448748 - INS 
 tpg|BK006949.2| 63047 + tpg|BK006949.2| 63712 - INS 
 tpg|BK006949.2| 223933 + tpg|BK006949.2| 223588 - INS 
 tpg|BK006949.2| 612972 + tpg|BK006949.2| 613628 - INS 
 tpg|BK006949.2| 730286 + tpg|BK006949.2| 730356 - INS 
 tpg|BK006949.2| 203413 + tpg|BK006949.2| 203026 - INS 
 tpg|BK006949.2| 444525 + tpg|BK006949.2| 444387 - INS 
 tpg|BK006949.2| 101677 + tpg|BK006949.2| 101180 - INS 
 tpg|BK006949.2| 398922 + tpg|BK006949.2| 398173 - INS 
 tpg|BK006949.2| 857706 + tpg|BK006949.2| 857194 - INS 
 tpg|BK006949.2| 828662 + tpg|BK006949.2| 828190 - INS 
 tpg|BK006949.2| 335722 + tpg|BK006949.2| 334961 - INS 
 tpg|BK006949.2| 328590 + tpg|BK006949.2| 329069 - INS 
 tpg|BK006949.2| 699196 + tpg|BK006949.2| 698982 - INS 
 tpg|BK006949.2| 410606 + tpg|BK006949.2| 410154 - INS 
 tpg|BK006949.2| 323615 + tpg|BK006949.2| 322951 - INS 
 tpg|BK006949.2| 663158 + tpg|BK006949.2| 662497 - INS 
 tpg|BK006949.2| 210714 + tpg|BK006949.2| 210817 - INS 
 tpg|BK006949.2| 307501 + tpg|BK006949.2| 306867 - INS 
 tpg|BK006949.2| 623577 + tpg|BK006949.2| 623214 - INS 
 tpg|BK006949.2| 605781 + tpg|BK006949.2| 605323 - INS 
 tpg|BK006949.2| 557490 + tpg|BK006949.2| 557360 - INS 
 tpg|BK006949.2| 892414 + tpg|BK006949.2| 893107 - INS 
 tpg|BK006949.2| 487991 + tpg|BK006949.2| 487775 - INS 
 tpg|BK006949.2| 532390 + tpg|BK006949.2| 532292 - INS 
 tpg|BK006949.2| 278335 + tpg|BK006949.2| 278145 - INS 
 tpg|BK006949.2| 316617 + tpg|BK006949.2| 316399 - INS 
 tpg|BK006949.2| 500968 + tpg|BK006949.2| 500808 - INS 
 tpg|BK006949.2| 242472 + tpg|BK006949.2| 242521 - INS 
 tpg|BK006949.2| 571586 + tpg|BK006949.2| 571180 - INS 
 tpg|BK006949.2| 156765 + tpg|BK006949.2| 156029 - INS 
 tpg|BK006949.2| 277708 + tpg|BK006949.2| 277186 - INS 
 tpg|BK006949.2| 537710 + tpg|BK006949.2| 538373 - INS 
 tpg|BK006949.2| 941344 + tpg|BK006949.2| 940626 - INS 
 tpg|BK006949.2| 923348 + tpg|BK006949.2| 923331 - INS 
 tpg|BK006949.2| 510729 + tpg|BK006949.2| 510546 - INS 
 tpg|BK006949.2| 261475 + tpg|BK006949.2| 260936 - INS 
 tpg|BK006949.2| 778300 + tpg|BK006949.2| 777608 - INS TC
 tpg|BK006949.2| 840194 + tpg|BK006949.2| 839900 - INS 
 tpg|BK006949.2| 255235 + tpg|BK006949.2| 255048 - INS 
 tpg|BK006949.2| 254307 + tpg|BK006949.2| 254063 - INS 
 tpg|BK006949.2| 147411 + tpg|BK006949.2| 147447 - INS 
 tpg|BK006949.2| 387478 + tpg|BK006949.2| 387640 - INS 
 tpg|BK006949.2| 417269 + tpg|BK006949.2| 416699 - INS 
 tpg|BK006949.2| 416549 + tpg|BK006949.2| 416199 - INS 
 tpg|BK006949.2| 632160 + tpg|BK006949.2| 632335 - INS 
 tpg|BK006949.2| 633123 + tpg|BK006949.2| 632783 - INS 
 tpg|BK006949.2| 641353 + tpg|BK006949.2| 640606 - INS 
 tpg|BK006949.2| 862275 + tpg|BK006949.2| 862429 - INS 
 tpg|BK006949.2| 97122 + tpg|BK006949.2| 96476 - INS 
 tpg|BK006949.2| 660799 + tpg|BK006949.2| 661450 - INS 
 tpg|BK006949.2| 341307 + tpg|BK006949.2| 340862 - INS 
 tpg|BK006949.2| 412487 + tpg|BK006949.2| 413170 - INS 
 tpg|BK006949.2| 866458 + tpg|BK006949.2| 865883 - INS 
 tpg|BK006949.2| 841204 + tpg|BK006949.2| 841427 - INS 
 tpg|BK006949.2| 411828 + tpg|BK006949.2| 411825 - INS 
 tpg|BK006949.2| 372609 + tpg|BK006949.2| 372555 - INS 
 tpg|BK006949.2| 869253 + tpg|BK006949.2| 869338 - INS 
 tpg|BK006949.2| 404123 + tpg|BK006949.2| 403681 - INS 
 tpg|BK006949.2| 160028 + tpg|BK006949.2| 159336 - INS 
 tpg|BK006949.2| 891228 + tpg|BK006949.2| 890973 - INS 
 tpg|BK006949.2| 622055 + tpg|BK006949.2| 621619 - INS 
 tpg|BK006949.2| 108292 + tpg|BK006949.2| 108757 - INS 
 tpg|BK006949.2| 443697 + tpg|BK006949.2| 443131 - INS 
 tpg|BK006949.2| 810844 + tpg|BK006949.2| 810486 - INS 
 tpg|BK006949.2| 26731 + tpg|BK006949.2| 26015 - INS 
 tpg|BK006949.2| 834243 + tpg|BK006949.2| 834840 - INS 
 tpg|BK006949.2| 746850 + tpg|BK006949.2| 746714 - INS 
 tpg|BK006949.2| 736664 + tpg|BK006949.2| 736211 - INS 
 tpg|BK006949.2| 595528 + tpg|BK006949.2| 595328 - INS 
 tpg|BK006949.2| 345811 + tpg|BK006949.2| 346089 - INS TAATGTTTGTG
 tpg|BK006949.2| 728163 + tpg|BK006949.2| 728171 - INS 
 tpg|BK006949.2| 726037 + tpg|BK006949.2| 726568 - INS 
 tpg|BK006949.2| 208459 + tpg|BK006949.2| 208109 - INS 
 tpg|BK006949.2| 169573 + tpg|BK006949.2| 169544 - INS 
 tpg|BK006949.2| 413968 + tpg|BK006949.2| 413621 - INS 
 tpg|BK006949.2| 431077 + tpg|BK006949.2| 430464 - INS 
 tpg|BK006949.2| 651016 + tpg|BK006949.2| 650325 - INS 
 tpg|BK006949.2| 308269 + tpg|BK006949.2| 307629 - INS 
 tpg|BK006949.2| 475030 + tpg|BK006949.2| 475325 - INS 
 tpg|BK006949.2| 116987 + tpg|BK006949.2| 116325 - INS 
 tpg|BK006949.2| 569335 + tpg|BK006949.2| 569961 - INS 
 tpg|BK006949.2| 236451 + tpg|BK006949.2| 236067 - INS 
 tpg|BK006949.2| 814837 + tpg|BK006949.2| 814782 - INS 
 tpg|BK006949.2| 368761 + tpg|BK006949.2| 368240 - INS 
 tpg|BK006949.2| 714518 + tpg|BK006949.2| 714812 - INS 
 tpg|BK006949.2| 524147 + tpg|BK006949.2| 523727 - INS 
 tpg|BK006949.2| 37062 + tpg|BK006949.2| 36412 - INS 
 tpg|BK006949.2| 499951 + tpg|BK006949.2| 499725 - INS 
 tpg|BK006949.2| 732500 + tpg|BK006949.2| 732737 - INS 
 tpg|BK006949.2| 495044 + tpg|BK006949.2| 494370 - INS 
 tpg|BK006949.2| 520184 + tpg|BK006949.2| 519566 - INS 
 tpg|BK006949.2| 365078 + tpg|BK006949.2| 364910 - INS 
 tpg|BK006949.2| 540041 + tpg|BK006949.2| 539807 - INS 
 tpg|BK006949.2| 400040 + tpg|BK006949.2| 399908 - INS 
 tpg|BK006949.2| 780277 + tpg|BK006949.2| 779808 - INS 
 tpg|BK006949.2| 544980 + tpg|BK006949.2| 544853 - INS 
 tpg|BK006949.2| 928786 + tpg|BK006949.2| 928263 - INS 
 tpg|BK006949.2| 145461 + tpg|BK006949.2| 144946 - INS 
 tpg|BK006949.2| 797350 + tpg|BK006949.2| 797979 - INS 
 tpg|BK006949.2| 685924 + tpg|BK006949.2| 686025 - INS 
 tpg|BK006949.2| 23691 + tpg|BK006949.2| 23328 - INS 
 tpg|BK006949.2| 864544 + tpg|BK006949.2| 864942 - INS 
 tpg|BK006949.2| 684877 + tpg|BK006949.2| 684527 - INS 
 tpg|BK006949.2| 908450 + tpg|BK006949.2| 908660 - INS 
 tpg|BK006949.2| 14846 + tpg|BK006949.2| 14969 - INS 
 tpg|BK006949.2| 602096 + tpg|BK006949.2| 601663 - INS 
 tpg|BK006949.2| 175563 + tpg|BK006949.2| 175496 - INS 
 tpg|BK006949.2| 507734 + tpg|BK006949.2| 508166 - INS 
 tpg|BK006949.2| 472478 + tpg|BK006949.2| 471887 - INS 
 tpg|BK006949.2| 422288 + tpg|BK006949.2| 421721 - INS 
 tpg|BK006949.2| 473380 + tpg|BK006949.2| 472717 - INS 
 tpg|BK006949.2| 941804 + tpg|BK006949.2| 941434 - INS 
 tpg|BK006949.2| 914059 + tpg|BK006949.2| 913498 - INS 
 tpg|BK006949.2| 588628 + tpg|BK006949.2| 588698 - INS 
 tpg|BK006949.2| 293552 + tpg|BK006949.2| 293812 - INS 
 tpg|BK006949.2| 942486 + tpg|BK006949.2| 942101 - INS 
 tpg|BK006949.2| 818865 + tpg|BK006949.2| 818776 - INS 
 tpg|BK006949.2| 449799 + tpg|BK006949.2| 450556 - INS 
 tpg|BK006949.2| 938418 + tpg|BK006949.2| 938389 - INS 
 tpg|BK006949.2| 82836 + tpg|BK006949.2| 82347 - INS 
 tpg|BK006949.2| 224505 + tpg|BK006949.2| 224310 - INS 
 tpg|BK006949.2| 665323 + tpg|BK006949.2| 664987 - INS 
 tpg|BK006949.2| 219271 + tpg|BK006949.2| 219119 - INS 
 tpg|BK006949.2| 913333 + tpg|BK006949.2| 912848 - INS 
 tpg|BK006949.2| 819672 + tpg|BK006949.2| 819666 - INS 
 tpg|BK006949.2| 375782 + tpg|BK006949.2| 375574 - INS 
 tpg|BK006949.2| 888934 + tpg|BK006949.2| 888884 - INS 
 tpg|BK006949.2| 38015 + tpg|BK006949.2| 37530 - INS 
 tpg|BK006949.2| 45684 + tpg|BK006949.2| 45068 - INS 
 tpg|BK006949.2| 757240 + tpg|BK006949.2| 757177 - INS 
 tpg|BK006949.2| 452662 + tpg|BK006949.2| 453089 - INS 
 tpg|BK006949.2| 702130 + tpg|BK006949.2| 701989 - INS 
 tpg|BK006949.2| 515162 + tpg|BK006949.2| 515337 - INS 
 tpg|BK006949.2| 312984 + tpg|BK006949.2| 313694 - INS 
 tpg|BK006949.2| 559857 + tpg|BK006949.2| 559954 - INS 
 tpg|BK006949.2| 838024 + tpg|BK006949.2| 837620 - INS 
 tpg|BK006949.2| 582220 + tpg|BK006949.2| 581713 - INS 
 tpg|BK006949.2| 577328 + tpg|BK006949.2| 577646 - INS 
 tpg|BK006949.2| 776292 + tpg|BK006949.2| 776367 - INS 
 tpg|BK006949.2| 228530 + tpg|BK006949.2| 227897 - INS 
 tpg|BK006949.2| 750726 + tpg|BK006949.2| 750922 - INS 
 tpg|BK006949.2| 408470 + tpg|BK006949.2| 407772 - INS 
 tpg|BK006949.2| 833267 + tpg|BK006949.2| 833926 - INS 
 tpg|BK006949.2| 255968 + tpg|BK006949.2| 255581 - INS 
 tpg|BK006949.2| 241746 + tpg|BK006949.2| 241596 - INS 
 tpg|BK006949.2| 354071 + tpg|BK006949.2| 353881 - INS 
 tpg|BK006949.2| 688932 + tpg|BK006949.2| 688727 - INS 
 tpg|BK006949.2| 826227 + tpg|BK006949.2| 826472 - INS 
 tpg|BK006949.2| 80237 + tpg|BK006949.2| 79544 - INS 
 tpg|BK006949.2| 593668 + tpg|BK006949.2| 593753 - INS 
 tpg|BK006949.2| 183271 + tpg|BK006949.2| 183391 - INS 
 tpg|BK006949.2| 625495 + tpg|BK006949.2| 625124 - INS 
 tpg|BK006949.2| 409167 + tpg|BK006949.2| 408675 - INS 
 tpg|BK006949.2| 924695 + tpg|BK006949.2| 924433 - INS 
 tpg|BK006949.2| 930154 + tpg|BK006949.2| 930578 - INS 
 tpg|BK006949.2| 751033 + tpg|BK006949.2| 751560 - INS 
 tpg|BK006949.2| 558708 + tpg|BK006949.2| 558863 - INS 
 tpg|BK006949.2| 170573 + tpg|BK006949.2| 169988 - INS 
 tpg|BK006949.2| 88136 + tpg|BK006949.2| 88074 - INS 
 tpg|BK006949.2| 93952 + tpg|BK006949.2| 93930 - INS 
 tpg|BK006949.2| 905956 + tpg|BK006949.2| 905949 - INS 
 tpg|BK006949.2| 858391 + tpg|BK006949.2| 857768 - INS 
 tpg|BK006949.2| 56405 + tpg|BK006949.2| 56373 - INS 
 tpg|BK006949.2| 304937 + tpg|BK006949.2| 305606 - INS 
 tpg|BK006949.2| 831706 + tpg|BK006949.2| 831299 - INS 
 tpg|BK006949.2| 925587 + tpg|BK006949.2| 925798 - INS 
 tpg|BK006949.2| 624052 + tpg|BK006949.2| 624719 - INS 
 tpg|BK006949.2| 70779 + tpg|BK006949.2| 70546 - INS 
 tpg|BK006949.2| 586299 + tpg|BK006949.2| 585547 - INS 
 tpg|BK006949.2| 762211 + tpg|BK006949.2| 762159 - INS 
 tpg|BK006949.2| 64734 + tpg|BK006949.2| 64922 - INS 
 tpg|BK006949.2| 509217 + tpg|BK006949.2| 509144 - INS 
 tpg|BK006949.2| 566528 + tpg|BK006949.2| 566285 - INS 
 tpg|BK006949.2| 877793 + tpg|BK006949.2| 877231 - INS 
 tpg|BK006949.2| 138513 + tpg|BK006949.2| 139085 - INS 
 tpg|BK006949.2| 140288 + tpg|BK006949.2| 140679 - INS 
 tpg|BK006949.2| 144124 + tpg|BK006949.2| 143668 - INS 
 tpg|BK006949.2| 663804 + tpg|BK006949.2| 663096 - INS 
 tpg|BK006949.2| 803394 + tpg|BK006949.2| 803013 - INS 
 tpg|BK006949.2| 286962 + tpg|BK006949.2| 287008 - INS 
 tpg|BK006949.2| 13764 + tpg|BK006949.2| 13174 - INS 
 tpg|BK006949.2| 844076 + tpg|BK006949.2| 843403 - INS 
 tpg|BK006949.2| 645689 + tpg|BK006949.2| 645965 - INS 
 tpg|BK006949.2| 683969 + tpg|BK006949.2| 683587 - INS 
 tpg|BK006949.2| 555339 + tpg|BK006949.2| 555412 - INS 
 tpg|BK006949.2| 909164 + tpg|BK006949.2| 909467 - INS 
 tpg|BK006949.2| 474027 + tpg|BK006949.2| 473382 - INS 
 tpg|BK006949.2| 918254 + tpg|BK006949.2| 917991 - INS 
 tpg|BK006949.2| 548017 + tpg|BK006949.2| 547608 - INS 
 tpg|BK006949.2| 266806 + tpg|BK006949.2| 267062 - INS 
 tpg|BK006949.2| 490756 + tpg|BK006949.2| 490705 - INS 
 tpg|BK006949.2| 690031 + tpg|BK006949.2| 690416 - INS 
 tpg|BK006949.2| 486897 + tpg|BK006949.2| 486944 - INS 
 tpg|BK006949.2| 29912 + tpg|BK006949.2| 29620 - INS 
 tpg|BK006949.2| 347533 + tpg|BK006949.2| 347029 - INS 
 tpg|BK006949.2| 820475 + tpg|BK006949.2| 820644 - INS 
 tpg|BK006949.2| 758727 + tpg|BK006949.2| 758254 - INS 
 tpg|BK006949.2| 274547 + tpg|BK006949.2| 274380 - INS 
 tpg|BK006949.2| 691981 + tpg|BK006949.2| 691892 - INS 
 tpg|BK006949.2| 162724 + tpg|BK006949.2| 163031 - INS 
 tpg|BK006949.2| 627591 + tpg|BK006949.2| 627523 - INS 
 tpg|BK006949.2| 240841 + tpg|BK006949.2| 240223 - INS 
 tpg|BK006949.2| 372022 + tpg|BK006949.2| 371793 - INS 
 tpg|BK006949.2| 44972 + tpg|BK006949.2| 44491 - INS 
 tpg|BK006949.2| 515832 + tpg|BK006949.2| 515939 - INS 
 tpg|BK006949.2| 416090 + tpg|BK006949.2| 415645 - INS 
 tpg|BK006949.2| 754914 + tpg|BK006949.2| 754486 - INS 
 tpg|BK006949.2| 576539 + tpg|BK006949.2| 576465 - INS 
 tpg|BK006949.2| 574457 + tpg|BK006949.2| 574453 - INS 
 tpg|BK006949.2| 850733 + tpg|BK006949.2| 850341 - INS 
 tpg|BK006949.2| 476930 + tpg|BK006949.2| 476719 - INS 
 tpg|BK006949.2| 72219 + tpg|BK006949.2| 71566 - INS 
 tpg|BK006949.2| 37734 + tpg|BK006949.2| 37086 - INS 
 tpg|BK006949.2| 119621 + tpg|BK006949.2| 118988 - INS 
 tpg|BK006949.2| 645046 + tpg|BK006949.2| 644806 - INS 
 tpg|BK006949.2| 249524 + tpg|BK006949.2| 249614 - INS 
 tpg|BK006949.2| 811286 + tpg|BK006949.2| 811240 - INS 
 tpg|BK006949.2| 724181 + tpg|BK006949.2| 724770 - INS 
 tpg|BK006949.2| 844537 + tpg|BK006949.2| 844006 - INS 
 tpg|BK006949.2| 741815 + tpg|BK006949.2| 741733 - INS 
 tpg|BK006949.2| 785391 + tpg|BK006949.2| 785719 - INS 
 tpg|BK006949.2| 315588 + tpg|BK006949.2| 315396 - INS 
 tpg|BK006949.2| 729248 + tpg|BK006949.2| 728599 - INS 
 tpg|BK006949.2| 342157 + tpg|BK006949.2| 342111 - INS 
 tpg|BK006949.2| 875249 + tpg|BK006949.2| 875393 - INS 
 tpg|BK006949.2| 181152 + tpg|BK006949.2| 181032 - INS 
 tpg|BK006948.2| 253164 + tpg|BK006948.2| 253735 - INS 
 tpg|BK006948.2| 96329 + tpg|BK006948.2| 97102 - INS 
 tpg|BK006948.2| 158175 + tpg|BK006948.2| 158828 - INS 
 tpg|BK006948.2| 1023107 + tpg|BK006948.2| 1022511 - INS 
 tpg|BK006948.2| 29073 + tpg|BK006948.2| 29829 - INS 
 tpg|BK006948.2| 1061644 + tpg|BK006948.2| 1061967 - INS 
 tpg|BK006948.2| 518599 + tpg|BK006948.2| 518161 - INS 
 tpg|BK006948.2| 638476 + tpg|BK006948.2| 637875 - INS 
 tpg|BK006948.2| 761473 + tpg|BK006948.2| 760961 - INS 
 tpg|BK006948.2| 797634 + tpg|BK006948.2| 796877 - INS 
 tpg|BK006948.2| 279363 + tpg|BK006948.2| 279353 - INS 
 tpg|BK006948.2| 352164 + tpg|BK006948.2| 351537 - INS 
 tpg|BK006948.2| 194290 + tpg|BK006948.2| 193661 - INS 
 tpg|BK006948.2| 208591 + tpg|BK006948.2| 209069 - INS 
 tpg|BK006948.2| 988356 + tpg|BK006948.2| 987870 - INS 
 tpg|BK006948.2| 410114 + tpg|BK006948.2| 409794 - INS 
 tpg|BK006948.2| 535434 + tpg|BK006948.2| 535346 - INS 
 tpg|BK006948.2| 305358 + tpg|BK006948.2| 305098 - INS 
 tpg|BK006948.2| 459030 + tpg|BK006948.2| 458979 - INS 
 tpg|BK006948.2| 1074091 + tpg|BK006948.2| 1073478 - INS 
 tpg|BK006948.2| 579990 + tpg|BK006948.2| 579255 - INS 
 tpg|BK006948.2| 162706 + tpg|BK006948.2| 162279 - INS 
 tpg|BK006948.2| 138355 + tpg|BK006948.2| 138900 - INS 
 tpg|BK006948.2| 146536 + tpg|BK006948.2| 146717 - INS 
 tpg|BK006948.2| 609235 + tpg|BK006948.2| 609621 - INS 
 tpg|BK006948.2| 514939 + tpg|BK006948.2| 515352 - INS 
 tpg|BK006948.2| 713379 + tpg|BK006948.2| 713369 - INS 
 tpg|BK006948.2| 890687 + tpg|BK006948.2| 891030 - INS 
 tpg|BK006948.2| 523367 + tpg|BK006948.2| 522803 - INS 
 tpg|BK006948.2| 646900 + tpg|BK006948.2| 646823 - INS 
 tpg|BK006948.2| 498839 + tpg|BK006948.2| 498084 - INS 
 tpg|BK006948.2| 488526 + tpg|BK006948.2| 487951 - INS 
 tpg|BK006948.2| 702478 + tpg|BK006948.2| 702010 - INS 
 tpg|BK006948.2| 451167 + tpg|BK006948.2| 450590 - INS 
 tpg|BK006948.2| 40979 + tpg|BK006948.2| 41298 - INS 
 tpg|BK006948.2| 794021 + tpg|BK006948.2| 793379 - INS 
 tpg|BK006948.2| 8971 + tpg|BK006948.2| 8539 - INS 
 tpg|BK006948.2| 688203 + tpg|BK006948.2| 688055 - INS 
 tpg|BK006948.2| 1006648 + tpg|BK006948.2| 1006751 - INS 
 tpg|BK006948.2| 1058374 + tpg|BK006948.2| 1059036 - INS 
 tpg|BK006948.2| 742652 + tpg|BK006948.2| 742825 - INS 
 tpg|BK006948.2| 377368 + tpg|BK006948.2| 376840 - INS 
 tpg|BK006948.2| 900905 + tpg|BK006948.2| 901068 - INS 
 tpg|BK006948.2| 907622 + tpg|BK006948.2| 907091 - INS 
 tpg|BK006948.2| 152490 + tpg|BK006948.2| 153078 - INS 
 tpg|BK006948.2| 57393 + tpg|BK006948.2| 57508 - INS 
 tpg|BK006948.2| 677094 + tpg|BK006948.2| 676903 - INS 
 tpg|BK006948.2| 46226 + tpg|BK006948.2| 45742 - INS 
 tpg|BK006948.2| 48522 + tpg|BK006948.2| 48970 - INS 
 tpg|BK006948.2| 460216 + tpg|BK006948.2| 460060 - INS 
 tpg|BK006948.2| 716394 + tpg|BK006948.2| 716967 - INS 
 tpg|BK006948.2| 25019 + tpg|BK006948.2| 24874 - INS 
 tpg|BK006948.2| 357282 + tpg|BK006948.2| 357547 - INS 
 tpg|BK006948.2| 772621 + tpg|BK006948.2| 773036 - INS 
 tpg|BK006948.2| 195773 + tpg|BK006948.2| 195201 - INS 
 tpg|BK006948.2| 334946 + tpg|BK006948.2| 334435 - INS 
 tpg|BK006948.2| 75844 + tpg|BK006948.2| 75707 - INS 
 tpg|BK006948.2| 276618 + tpg|BK006948.2| 276169 - INS 
 tpg|BK006948.2| 81344 + tpg|BK006948.2| 80951 - INS 
 tpg|BK006948.2| 225025 + tpg|BK006948.2| 224688 - INS 
 tpg|BK006948.2| 829904 + tpg|BK006948.2| 830577 - INS 
 tpg|BK006948.2| 938100 + tpg|BK006948.2| 937574 - INS 
 tpg|BK006948.2| 652558 + tpg|BK006948.2| 653168 - INS 
 tpg|BK006948.2| 562816 + tpg|BK006948.2| 562181 - INS 
 tpg|BK006948.2| 898412 + tpg|BK006948.2| 898584 - INS 
 tpg|BK006948.2| 441443 + tpg|BK006948.2| 441720 - INS 
 tpg|BK006948.2| 712460 + tpg|BK006948.2| 711952 - INS 
 tpg|BK006948.2| 205747 + tpg|BK006948.2| 205846 - INS 
 tpg|BK006948.2| 834267 + tpg|BK006948.2| 833604 - INS 
 tpg|BK006948.2| 737584 + tpg|BK006948.2| 738330 - INS 
 tpg|BK006948.2| 312040 + tpg|BK006948.2| 311945 - INS 
 tpg|BK006948.2| 425350 + tpg|BK006948.2| 425548 - INS 
 tpg|BK006948.2| 6174 + tpg|BK006948.2| 6532 - INS 
 tpg|BK006948.2| 494732 + tpg|BK006948.2| 494200 - INS 
 tpg|BK006948.2| 744450 + tpg|BK006948.2| 744190 - INS 
 tpg|BK006948.2| 955078 + tpg|BK006948.2| 955043 - INS 
 tpg|BK006948.2| 553358 + tpg|BK006948.2| 553249 - INS 
 tpg|BK006948.2| 636625 + tpg|BK006948.2| 636885 - INS 
 tpg|BK006948.2| 462339 + tpg|BK006948.2| 461865 - INS 
 tpg|BK006948.2| 897198 + tpg|BK006948.2| 897051 - INS 
 tpg|BK006948.2| 578233 + tpg|BK006948.2| 577591 - INS 
 tpg|BK006948.2| 689373 + tpg|BK006948.2| 688967 - INS 
 tpg|BK006948.2| 440718 + tpg|BK006948.2| 441088 - INS 
 tpg|BK006948.2| 417591 + tpg|BK006948.2| 417637 - INS 
 tpg|BK006948.2| 814728 + tpg|BK006948.2| 814078 - INS 
 tpg|BK006948.2| 819341 + tpg|BK006948.2| 819233 - INS 
 tpg|BK006948.2| 872387 + tpg|BK006948.2| 873111 - INS 
 ref|NC_001224| 17189 + ref|NC_001224| 16961 - INS 
 tpg|BK006948.2| 954364 + tpg|BK006948.2| 954152 - INS 
 tpg|BK006948.2| 210347 + tpg|BK006948.2| 209868 - INS 
 tpg|BK006948.2| 457410 + tpg|BK006948.2| 456813 - INS 
 tpg|BK006948.2| 391963 + tpg|BK006948.2| 391437 - INS 
 tpg|BK006948.2| 362103 + tpg|BK006948.2| 361809 - INS 
 tpg|BK006948.2| 1002316 + tpg|BK006948.2| 1002241 - INS 
 tpg|BK006948.2| 906819 + tpg|BK006948.2| 906548 - INS 
 tpg|BK006948.2| 272466 + tpg|BK006948.2| 271704 - INS 
 tpg|BK006948.2| 264590 + tpg|BK006948.2| 264399 - INS 
 tpg|BK006948.2| 213271 + tpg|BK006948.2| 212716 - INS 
 tpg|BK006948.2| 1069147 + tpg|BK006948.2| 1068429 - INS 
 tpg|BK006948.2| 836361 + tpg|BK006948.2| 836020 - INS 
 tpg|BK006948.2| 546091 + tpg|BK006948.2| 546004 - INS 
 tpg|BK006948.2| 1030340 + tpg|BK006948.2| 1030387 - INS 
 tpg|BK006948.2| 883257 + tpg|BK006948.2| 883119 - INS 
 tpg|BK006948.2| 559818 + tpg|BK006948.2| 559091 - INS 
 tpg|BK006948.2| 473171 + tpg|BK006948.2| 473221 - INS 
 tpg|BK006948.2| 306303 + tpg|BK006948.2| 306420 - INS 
 tpg|BK006948.2| 502284 + tpg|BK006948.2| 502703 - INS 
 tpg|BK006948.2| 544431 + tpg|BK006948.2| 544285 - INS 
 tpg|BK006948.2| 668929 + tpg|BK006948.2| 668539 - INS 
 tpg|BK006948.2| 669462 + tpg|BK006948.2| 669091 - INS 
 tpg|BK006948.2| 468738 + tpg|BK006948.2| 469423 - INS 
 tpg|BK006948.2| 720205 + tpg|BK006948.2| 719491 - INS 
 tpg|BK006948.2| 655305 + tpg|BK006948.2| 654911 - INS 
 tpg|BK006948.2| 692084 + tpg|BK006948.2| 691856 - INS 
 tpg|BK006948.2| 230569 + tpg|BK006948.2| 230509 - INS 
 tpg|BK006948.2| 448362 + tpg|BK006948.2| 448398 - INS 
 tpg|BK006948.2| 747827 + tpg|BK006948.2| 748546 - INS 
 tpg|BK006948.2| 92472 + tpg|BK006948.2| 92774 - INS 
 tpg|BK006948.2| 788196 + tpg|BK006948.2| 787901 - INS 
 tpg|BK006948.2| 792428 + tpg|BK006948.2| 791810 - INS 
 tpg|BK006948.2| 1027576 + tpg|BK006948.2| 1027238 - INS 
 tpg|BK006948.2| 71087 + tpg|BK006948.2| 70535 - INS 
 tpg|BK006948.2| 893860 + tpg|BK006948.2| 893516 - INS 
 tpg|BK006948.2| 248959 + tpg|BK006948.2| 248235 - INS 
 tpg|BK006948.2| 928613 + tpg|BK006948.2| 928218 - INS 
 tpg|BK006948.2| 690065 + tpg|BK006948.2| 689826 - INS 
 tpg|BK006948.2| 724391 + tpg|BK006948.2| 725106 - INS 
 tpg|BK006948.2| 521687 + tpg|BK006948.2| 522133 - INS 
 tpg|BK006948.2| 933225 + tpg|BK006948.2| 932643 - INS 
 tpg|BK006948.2| 726022 + tpg|BK006948.2| 725878 - INS 
 tpg|BK006948.2| 314617 + tpg|BK006948.2| 314885 - INS 
 tpg|BK006948.2| 104856 + tpg|BK006948.2| 105054 - INS 
 tpg|BK006948.2| 389042 + tpg|BK006948.2| 389565 - INS 
 tpg|BK006948.2| 427028 + tpg|BK006948.2| 427176 - INS 
 tpg|BK006948.2| 626126 + tpg|BK006948.2| 626663 - INS 
 tpg|BK006939.2| 504118 + tpg|BK006939.2| 504157 - INS 
 tpg|BK006948.2| 408688 + tpg|BK006948.2| 409338 - INS 
 tpg|BK006948.2| 380766 + tpg|BK006948.2| 381132 - INS 
 tpg|BK006948.2| 333445 + tpg|BK006948.2| 333842 - INS 
 tpg|BK006948.2| 317970 + tpg|BK006948.2| 318500 - INS 
 tpg|BK006948.2| 984660 + tpg|BK006948.2| 984787 - INS 
 tpg|BK006948.2| 583440 + tpg|BK006948.2| 582757 - INS 
 tpg|BK006948.2| 1044171 + tpg|BK006948.2| 1043400 - INS 
 tpg|BK006948.2| 173121 + tpg|BK006948.2| 173667 - INS 
 tpg|BK006948.2| 4095 + tpg|BK006948.2| 4081 - INS 
 tpg|BK006939.2| 322219 + tpg|BK006939.2| 321509 - INS 
 tpg|BK006939.2| 34338 + tpg|BK006939.2| 34026 - INS 
 tpg|BK006948.2| 43001 + tpg|BK006948.2| 42468 - INS 
 tpg|BK006948.2| 296298 + tpg|BK006948.2| 296787 - INS 
 tpg|BK006939.2| 400860 + tpg|BK006939.2| 400425 - INS 
 tpg|BK006948.2| 165064 + tpg|BK006948.2| 165516 - INS 
 tpg|BK006948.2| 107248 + tpg|BK006948.2| 106565 - INS 
 tpg|BK006948.2| 895033 + tpg|BK006948.2| 895377 - INS 
 tpg|BK006948.2| 403858 + tpg|BK006948.2| 404343 - INS 
 tpg|BK006948.2| 182157 + tpg|BK006948.2| 181632 - INS 
 tpg|BK006948.2| 424013 + tpg|BK006948.2| 424261 - INS 
 tpg|BK006948.2| 536147 + tpg|BK006948.2| 536894 - INS 
 tpg|BK006939.2| 122742 + tpg|BK006939.2| 123205 - INS 
 tpg|BK006948.2| 495671 + tpg|BK006948.2| 495702 - INS 
 tpg|BK006939.2| 42873 + tpg|BK006939.2| 42746 - INS 
 tpg|BK006948.2| 202606 + tpg|BK006948.2| 203036 - INS 
 tpg|BK006939.2| 126512 + tpg|BK006939.2| 126424 - INS 
 tpg|BK006939.2| 59815 + tpg|BK006939.2| 59428 - INS 
 tpg|BK006948.2| 215034 + tpg|BK006948.2| 215226 - INS 
 tpg|BK006939.2| 279701 + tpg|BK006939.2| 279484 - INS 
 tpg|BK006948.2| 64387 + tpg|BK006948.2| 64526 - INS 
 tpg|BK006948.2| 750527 + tpg|BK006948.2| 750589 - INS 
 tpg|BK006939.2| 462300 + tpg|BK006939.2| 463009 - INS 
 tpg|BK006948.2| 257864 + tpg|BK006948.2| 257944 - INS 
 tpg|BK006939.2| 475492 + tpg|BK006939.2| 474825 - INS 
 tpg|BK006948.2| 156162 + tpg|BK006948.2| 156184 - INS 
 tpg|BK006948.2| 888982 + tpg|BK006948.2| 888412 - INS 
 tpg|BK006948.2| 269987 + tpg|BK006948.2| 269799 - INS 
 tpg|BK006948.2| 990794 + tpg|BK006948.2| 990470 - INS 
 tpg|BK006948.2| 607906 + tpg|BK006948.2| 608644 - INS 
 tpg|BK006948.2| 613781 + tpg|BK006948.2| 614218 - INS 
 tpg|BK006939.2| 543039 + tpg|BK006939.2| 543141 - INS 
 tpg|BK006948.2| 1067257 + tpg|BK006948.2| 1066760 - INS 
 tpg|BK006939.2| 461614 + tpg|BK006939.2| 460953 - INS 
 tpg|BK006948.2| 1028194 + tpg|BK006948.2| 1028777 - INS 
 tpg|BK006948.2| 378120 + tpg|BK006948.2| 378004 - INS 
 tpg|BK006939.2| 411564 + tpg|BK006939.2| 411258 - INS 
 tpg|BK006948.2| 381596 + tpg|BK006948.2| 381803 - INS 
 tpg|BK006939.2| 415767 + tpg|BK006939.2| 416205 - INS 
 tpg|BK006948.2| 1034714 + tpg|BK006948.2| 1033965 - INS 
 tpg|BK006939.2| 418256 + tpg|BK006939.2| 418263 - INS 
 tpg|BK006948.2| 127946 + tpg|BK006948.2| 127998 - INS 
 tpg|BK006939.2| 526108 + tpg|BK006939.2| 526653 - INS 
 tpg|BK006948.2| 763363 + tpg|BK006948.2| 762791 - INS 
 tpg|BK006948.2| 108936 + tpg|BK006948.2| 108456 - INS 
 tpg|BK006939.2| 457389 + tpg|BK006939.2| 456853 - INS 
 tpg|BK006948.2| 38766 + tpg|BK006948.2| 38647 - INS 
 tpg|BK006939.2| 222936 + tpg|BK006939.2| 222650 - INS 
 tpg|BK006939.2| 41213 + tpg|BK006939.2| 41105 - INS 
 tpg|BK006939.2| 209936 + tpg|BK006939.2| 209258 - INS 
 tpg|BK006939.2| 329719 + tpg|BK006939.2| 328974 - INS 
 tpg|BK006948.2| 777247 + tpg|BK006948.2| 776802 - INS 
 tpg|BK006939.2| 70406 + tpg|BK006939.2| 70484 - INS 
 tpg|BK006948.2| 144064 + tpg|BK006948.2| 143829 - INS 
 tpg|BK006948.2| 741339 + tpg|BK006948.2| 741803 - INS 
 tpg|BK006948.2| 861813 + tpg|BK006948.2| 861770 - INS 
 tpg|BK006939.2| 240835 + tpg|BK006939.2| 240372 - INS 
 tpg|BK006948.2| 292591 + tpg|BK006948.2| 292874 - INS 
 tpg|BK006939.2| 117829 + tpg|BK006939.2| 117708 - INS 
 tpg|BK006948.2| 289019 + tpg|BK006948.2| 289291 - INS 
 tpg|BK006948.2| 612863 + tpg|BK006948.2| 612264 - INS 
 tpg|BK006939.2| 79223 + tpg|BK006939.2| 79689 - INS 
 tpg|BK006948.2| 530223 + tpg|BK006948.2| 530790 - INS AAG
 tpg|BK006948.2| 900158 + tpg|BK006948.2| 900261 - INS 
 tpg|BK006939.2| 376891 + tpg|BK006939.2| 376332 - INS 
 tpg|BK006948.2| 170938 + tpg|BK006948.2| 170763 - INS 
 tpg|BK006948.2| 524297 + tpg|BK006948.2| 523822 - INS 
 tpg|BK006939.2| 372335 + tpg|BK006939.2| 372931 - INS 
 tpg|BK006948.2| 164583 + tpg|BK006948.2| 163821 - INS 
 tpg|BK006948.2| 841700 + tpg|BK006948.2| 841153 - INS 
 tpg|BK006939.2| 269708 + tpg|BK006939.2| 269265 - INS 
 tpg|BK006948.2| 242256 + tpg|BK006948.2| 241945 - INS 
 tpg|BK006939.2| 187403 + tpg|BK006939.2| 187372 - INS 
 tpg|BK006939.2| 551973 + tpg|BK006939.2| 552718 - INS 
 tpg|BK006948.2| 181215 + tpg|BK006948.2| 180941 - INS 
 tpg|BK006948.2| 993714 + tpg|BK006948.2| 994384 - INS 
 tpg|BK006939.2| 433193 + tpg|BK006939.2| 433668 - INS 
 tpg|BK006948.2| 480202 + tpg|BK006948.2| 480150 - INS 
 tpg|BK006948.2| 32002 + tpg|BK006948.2| 31785 - INS 
 tpg|BK006939.2| 145112 + tpg|BK006939.2| 144749 - INS 
 tpg|BK006939.2| 200074 + tpg|BK006939.2| 199707 - INS 
 tpg|BK006939.2| 540417 + tpg|BK006939.2| 539972 - INS 
 tpg|BK006948.2| 402393 + tpg|BK006948.2| 402101 - INS 
 tpg|BK006939.2| 52250 + tpg|BK006939.2| 52059 - INS 
 tpg|BK006948.2| 1036017 + tpg|BK006948.2| 1036612 - INS 
 tpg|BK006939.2| 389249 + tpg|BK006939.2| 388910 - INS 
 tpg|BK006948.2| 1016418 + tpg|BK006948.2| 1016409 - INS 
 tpg|BK006939.2| 133745 + tpg|BK006939.2| 134285 - INS 
 tpg|BK006948.2| 718654 + tpg|BK006948.2| 718205 - INS 
 tpg|BK006939.2| 350968 + tpg|BK006939.2| 350632 - INS 
 tpg|BK006948.2| 918895 + tpg|BK006948.2| 918487 - INS 
 tpg|BK006939.2| 484945 + tpg|BK006939.2| 485075 - INS 
 tpg|BK006948.2| 1026746 + tpg|BK006948.2| 1026210 - INS 
 tpg|BK006939.2| 27709 + tpg|BK006939.2| 27363 - INS 
 tpg|BK006948.2| 384554 + tpg|BK006948.2| 384542 - INS 
 tpg|BK006948.2| 909188 + tpg|BK006948.2| 909376 - INS 
 tpg|BK006939.2| 489150 + tpg|BK006939.2| 489546 - INS 
 tpg|BK006948.2| 184823 + tpg|BK006948.2| 184451 - INS 
 tpg|BK006939.2| 160664 + tpg|BK006939.2| 160420 - INS 
 tpg|BK006948.2| 768114 + tpg|BK006948.2| 767488 - INS 
 tpg|BK006939.2| 507341 + tpg|BK006939.2| 507571 - INS 
 tpg|BK006939.2| 522387 + tpg|BK006939.2| 522819 - INS 
 tpg|BK006939.2| 479532 + tpg|BK006939.2| 480229 - INS 
 tpg|BK006948.2| 943217 + tpg|BK006948.2| 943129 - INS 
 tpg|BK006939.2| 510051 + tpg|BK006939.2| 510553 - INS 
 tpg|BK006948.2| 940352 + tpg|BK006948.2| 939830 - INS 
 tpg|BK006948.2| 903218 + tpg|BK006948.2| 903756 - INS 
 tpg|BK006939.2| 184087 + tpg|BK006939.2| 183691 - INS 
 tpg|BK006948.2| 916857 + tpg|BK006948.2| 917422 - INS 
 tpg|BK006939.2| 99232 + tpg|BK006939.2| 98947 - INS 
 tpg|BK006948.2| 1055063 + tpg|BK006948.2| 1055772 - INS 
 tpg|BK006948.2| 513258 + tpg|BK006948.2| 512552 - INS 
 tpg|BK006939.2| 564335 + tpg|BK006939.2| 564109 - INS 
 tpg|BK006948.2| 453697 + tpg|BK006948.2| 453556 - INS 
 tpg|BK006939.2| 331838 + tpg|BK006939.2| 331766 - INS 
 tpg|BK006948.2| 1065126 + tpg|BK006948.2| 1064565 - INS 
 tpg|BK006939.2| 349366 + tpg|BK006939.2| 349936 - INS 
 tpg|BK006948.2| 379824 + tpg|BK006948.2| 379801 - INS 
 tpg|BK006948.2| 445250 + tpg|BK006948.2| 444619 - INS 
 tpg|BK006939.2| 102814 + tpg|BK006939.2| 103185 - INS 
 tpg|BK006948.2| 434741 + tpg|BK006948.2| 434014 - INS 
 tpg|BK006939.2| 223819 + tpg|BK006939.2| 223690 - INS 
 tpg|BK006939.2| 453599 + tpg|BK006939.2| 452971 - INS 
 tpg|BK006939.2| 29347 + tpg|BK006939.2| 28666 - INS 
 tpg|BK006948.2| 481591 + tpg|BK006948.2| 481237 - INS 
 tpg|BK006948.2| 220581 + tpg|BK006948.2| 221070 - INS 
 tpg|BK006948.2| 211421 + tpg|BK006948.2| 211080 - INS 
 tpg|BK006948.2| 44219 + tpg|BK006948.2| 43807 - INS 
 tpg|BK006939.2| 161475 + tpg|BK006939.2| 162120 - INS 
 tpg|BK006948.2| 1051238 + tpg|BK006948.2| 1050738 - INS 
 tpg|BK006948.2| 217080 + tpg|BK006948.2| 217096 - INS 
 tpg|BK006939.2| 197337 + tpg|BK006939.2| 196607 - INS 
 tpg|BK006948.2| 443027 + tpg|BK006948.2| 442499 - INS 
 tpg|BK006939.2| 192218 + tpg|BK006939.2| 191915 - INS 
 tpg|BK006939.2| 57373 + tpg|BK006939.2| 57720 - INS 
 tpg|BK006939.2| 353977 + tpg|BK006939.2| 353277 - INS 
 tpg|BK006948.2| 273327 + tpg|BK006948.2| 273600 - INS 
 tpg|BK006939.2| 35780 + tpg|BK006939.2| 35599 - INS 
 tpg|BK006948.2| 1038276 + tpg|BK006948.2| 1037655 - INS 
 tpg|BK006939.2| 30727 + tpg|BK006939.2| 31266 - INS 
 tpg|BK006948.2| 228126 + tpg|BK006948.2| 228432 - INS 
 tpg|BK006948.2| 392828 + tpg|BK006948.2| 392454 - INS 
 tpg|BK006939.2| 402216 + tpg|BK006939.2| 402050 - INS 
 tpg|BK006948.2| 142918 + tpg|BK006948.2| 142250 - INS 
 tpg|BK006939.2| 90932 + tpg|BK006939.2| 91656 - INS 
 tpg|BK006948.2| 818100 + tpg|BK006948.2| 817594 - INS 
 tpg|BK006948.2| 321622 + tpg|BK006948.2| 321595 - INS 
 tpg|BK006948.2| 317069 + tpg|BK006948.2| 316776 - INS 
 tpg|BK006948.2| 299540 + tpg|BK006948.2| 299450 - INS 
 tpg|BK006948.2| 865696 + tpg|BK006948.2| 865895 - INS 
 tpg|BK006948.2| 78781 + tpg|BK006948.2| 78942 - INS 
 tpg|BK006948.2| 998004 + tpg|BK006948.2| 998108 - INS 
 tpg|BK006948.2| 879434 + tpg|BK006948.2| 878842 - INS 
 tpg|BK006939.2| 237733 + tpg|BK006939.2| 237840 - INS 
 tpg|BK006948.2| 627037 + tpg|BK006948.2| 627096 - INS 
 tpg|BK006939.2| 336835 + tpg|BK006939.2| 336119 - INS 
 tpg|BK006948.2| 192617 + tpg|BK006948.2| 192987 - INS 
 tpg|BK006939.2| 513453 + tpg|BK006939.2| 513399 - INS 
 tpg|BK006948.2| 967531 + tpg|BK006948.2| 967112 - INS 
 tpg|BK006939.2| 145533 + tpg|BK006939.2| 146008 - INS 
 tpg|BK006948.2| 656384 + tpg|BK006948.2| 656574 - INS 
 tpg|BK006948.2| 663448 + tpg|BK006948.2| 662765 - INS 
 tpg|BK006939.2| 198402 + tpg|BK006939.2| 198486 - INS 
 tpg|BK006948.2| 573430 + tpg|BK006948.2| 572673 - INS 
 tpg|BK006948.2| 1074509 + tpg|BK006948.2| 1074315 - INS 
 tpg|BK006939.2| 534670 + tpg|BK006939.2| 534622 - INS 
 tpg|BK006948.2| 199864 + tpg|BK006948.2| 200532 - INS 
 tpg|BK006939.2| 337462 + tpg|BK006939.2| 337652 - INS 
 tpg|BK006948.2| 348654 + tpg|BK006948.2| 348310 - INS 
 tpg|BK006939.2| 567939 + tpg|BK006939.2| 567659 - INS 
 tpg|BK006948.2| 801744 + tpg|BK006948.2| 801609 - INS 
 tpg|BK006948.2| 352971 + tpg|BK006948.2| 352238 - INS 
 tpg|BK006939.2| 265335 + tpg|BK006939.2| 265016 - INS 
 tpg|BK006948.2| 601353 + tpg|BK006948.2| 600837 - INS 
 tpg|BK006939.2| 237038 + tpg|BK006939.2| 236697 - INS 
 tpg|BK006948.2| 171682 + tpg|BK006948.2| 171852 - INS 
 tpg|BK006948.2| 683232 + tpg|BK006948.2| 682740 - INS 
 tpg|BK006948.2| 371191 + tpg|BK006948.2| 371862 - INS 
 tpg|BK006948.2| 585011 + tpg|BK006948.2| 585440 - INS 
 tpg|BK006939.2| 405860 + tpg|BK006939.2| 405278 - INS 
 tpg|BK006948.2| 416739 + tpg|BK006948.2| 416096 - INS 
 tpg|BK006939.2| 201941 + tpg|BK006939.2| 201668 - INS 
 tpg|BK006948.2| 65679 + tpg|BK006948.2| 65228 - INS 
 tpg|BK006948.2| 490439 + tpg|BK006948.2| 490163 - INS 
 tpg|BK006939.2| 378463 + tpg|BK006939.2| 378297 - INS 
 tpg|BK006948.2| 115153 + tpg|BK006948.2| 115459 - INS 
 tpg|BK006948.2| 1045456 + tpg|BK006948.2| 1045093 - INS 
 tpg|BK006948.2| 774217 + tpg|BK006948.2| 774766 - INS 
 tpg|BK006939.2| 278643 + tpg|BK006939.2| 278517 - INS 
 tpg|BK006948.2| 1049516 + tpg|BK006948.2| 1049435 - INS 
 tpg|BK006939.2| 424485 + tpg|BK006939.2| 424616 - INS 
 tpg|BK006948.2| 131994 + tpg|BK006948.2| 131406 - INS 
 tpg|BK006948.2| 1039268 + tpg|BK006948.2| 1038696 - INS 
 tpg|BK006939.2| 426109 + tpg|BK006939.2| 426425 - INS 
 tpg|BK006948.2| 839356 + tpg|BK006948.2| 839035 - INS 
 tpg|BK006939.2| 554521 + tpg|BK006939.2| 554201 - INS 
 tpg|BK006939.2| 32556 + tpg|BK006939.2| 32139 - INS 
 tpg|BK006948.2| 151463 + tpg|BK006948.2| 150928 - INS 
 tpg|BK006948.2| 307456 + tpg|BK006948.2| 307518 - INS 
 tpg|BK006939.2| 15260 + tpg|BK006939.2| 14621 - INS 
 tpg|BK006948.2| 368526 + tpg|BK006948.2| 367924 - INS 
 tpg|BK006939.2| 386153 + tpg|BK006939.2| 386138 - INS 
 tpg|BK006948.2| 740149 + tpg|BK006948.2| 740062 - INS 
 tpg|BK006939.2| 361709 + tpg|BK006939.2| 361888 - INS 
 tpg|BK006939.2| 541253 + tpg|BK006939.2| 542000 - INS 
 tpg|BK006939.2| 230221 + tpg|BK006939.2| 230054 - INS 
 tpg|BK006948.2| 337694 + tpg|BK006948.2| 337622 - INS 
 tpg|BK006939.2| 119594 + tpg|BK006939.2| 119482 - INS 
 tpg|BK006939.2| 359518 + tpg|BK006939.2| 358777 - INS 
 tpg|BK006948.2| 858151 + tpg|BK006948.2| 858496 - INS 
 tpg|BK006939.2| 431021 + tpg|BK006939.2| 430660 - INS 
 tpg|BK006948.2| 915960 + tpg|BK006948.2| 915920 - INS 
 tpg|BK006939.2| 67868 + tpg|BK006939.2| 67866 - INS 
 tpg|BK006948.2| 243715 + tpg|BK006948.2| 244282 - INS 
 tpg|BK006939.2| 490708 + tpg|BK006939.2| 490255 - INS 
 tpg|BK006948.2| 878093 + tpg|BK006948.2| 877622 - INS 
 ref|NC_001224| 16560 + ref|NC_001224| 16354 - INS 
 tpg|BK006939.2| 481267 + tpg|BK006939.2| 481818 - INS 
 tpg|BK006948.2| 13951 + tpg|BK006948.2| 13471 - INS 
 tpg|BK006939.2| 505589 + tpg|BK006939.2| 505849 - INS 
 tpg|BK006948.2| 699122 + tpg|BK006948.2| 698762 - INS 
 tpg|BK006939.2| 97852 + tpg|BK006939.2| 98227 - INS 
 tpg|BK006948.2| 422864 + tpg|BK006948.2| 423201 - INS 
 tpg|BK006939.2| 459175 + tpg|BK006939.2| 458891 - INS 
 tpg|BK006948.2| 541976 + tpg|BK006948.2| 542705 - INS 
 tpg|BK006939.2| 529329 + tpg|BK006939.2| 528595 - INS 
 tpg|BK006939.2| 544985 + tpg|BK006939.2| 545224 - INS 
 tpg|BK006939.2| 569053 + tpg|BK006939.2| 569684 - INS 
 tpg|BK006939.2| 427646 + tpg|BK006939.2| 427369 - INS 
 tpg|BK006939.2| 310802 + tpg|BK006939.2| 310314 - INS 
 tpg|BK006939.2| 143682 + tpg|BK006939.2| 143963 - INS 
 tpg|BK006948.2| 482759 + tpg|BK006948.2| 483133 - INS 
 tpg|BK006939.2| 267456 + tpg|BK006939.2| 267326 - INS 
 tpg|BK006939.2| 76188 + tpg|BK006939.2| 75846 - INS 
 tpg|BK006948.2| 88950 + tpg|BK006948.2| 88360 - INS 
 tpg|BK006939.2| 157033 + tpg|BK006939.2| 156337 - INS 
 tpg|BK006948.2| 213837 + tpg|BK006948.2| 214163 - INS 
 tpg|BK006939.2| 244807 + tpg|BK006939.2| 244563 - INS 
 tpg|BK006948.2| 445850 + tpg|BK006948.2| 445310 - INS 
 tpg|BK006939.2| 50817 + tpg|BK006939.2| 51402 - INS 
 tpg|BK006948.2| 589249 + tpg|BK006948.2| 588650 - INS 
 tpg|BK006939.2| 549320 + tpg|BK006939.2| 549226 - INS 
 tpg|BK006939.2| 516768 + tpg|BK006939.2| 516006 - INS 
 tpg|BK006948.2| 403080 + tpg|BK006948.2| 402982 - INS 
 tpg|BK006939.2| 174512 + tpg|BK006939.2| 174916 - INS 
 tpg|BK006948.2| 421621 + tpg|BK006948.2| 422316 - INS 
 tpg|BK006939.2| 473769 + tpg|BK006939.2| 473008 - INS 
 tpg|BK006939.2| 207325 + tpg|BK006939.2| 207228 - INS 
 tpg|BK006948.2| 397241 + tpg|BK006948.2| 397478 - INS 
 tpg|BK006948.2| 360524 + tpg|BK006948.2| 359841 - INS 
 tpg|BK006939.2| 47289 + tpg|BK006939.2| 47858 - INS 
 tpg|BK006948.2| 354302 + tpg|BK006948.2| 353743 - INS 
 tpg|BK006948.2| 267731 + tpg|BK006948.2| 268217 - INS 
 tpg|BK006939.2| 482984 + tpg|BK006939.2| 482624 - INS GAAAG
 tpg|BK006939.2| 53752 + tpg|BK006939.2| 53454 - INS 
 tpg|BK006948.2| 290282 + tpg|BK006948.2| 290742 - INS 
 tpg|BK006939.2| 369113 + tpg|BK006939.2| 368911 - INS 
 tpg|BK006939.2| 483869 + tpg|BK006939.2| 483453 - INS 
 tpg|BK006948.2| 2789 + tpg|BK006948.2| 2633 - INS 
 tpg|BK006939.2| 281108 + tpg|BK006939.2| 280926 - INS 
 tpg|BK006939.2| 340429 + tpg|BK006939.2| 339735 - INS 
 tpg|BK006939.2| 241868 + tpg|BK006939.2| 241727 - INS 
 tpg|BK006939.2| 330276 + tpg|BK006939.2| 329890 - INS 
 tpg|BK006948.2| 102993 + tpg|BK006948.2| 103512 - INS 
 tpg|BK006948.2| 849472 + tpg|BK006948.2| 849052 - INS 
 tpg|BK006939.2| 129930 + tpg|BK006939.2| 129834 - INS 
 tpg|BK006948.2| 628380 + tpg|BK006948.2| 627973 - INS 
 tpg|BK006939.2| 157765 + tpg|BK006939.2| 158394 - INS 
 tpg|BK006948.2| 250858 + tpg|BK006948.2| 251073 - INS 
 tpg|BK006948.2| 192046 + tpg|BK006948.2| 191750 - INS 
 tpg|BK006939.2| 325513 + tpg|BK006939.2| 325176 - INS 
 tpg|BK006948.2| 827130 + tpg|BK006948.2| 826841 - INS 
 tpg|BK006939.2| 501904 + tpg|BK006939.2| 501734 - INS 
 tpg|BK006939.2| 72980 + tpg|BK006939.2| 72432 - INS 
 tpg|BK006939.2| 550765 + tpg|BK006939.2| 550441 - INS 
 tpg|BK006939.2| 215343 + tpg|BK006939.2| 214614 - INS 
 tpg|BK006939.2| 63125 + tpg|BK006939.2| 63693 - INS 
 tpg|BK006948.2| 651611 + tpg|BK006948.2| 651070 - INS 
 tpg|BK006948.2| 7510 + tpg|BK006948.2| 8021 - INS 
 tpg|BK006939.2| 291901 + tpg|BK006939.2| 292058 - INS 
 tpg|BK006939.2| 212665 + tpg|BK006939.2| 212089 - INS 
 tpg|BK006948.2| 285704 + tpg|BK006948.2| 285142 - INS 
 tpg|BK006948.2| 826013 + tpg|BK006948.2| 826207 - INS 
 tpg|BK006939.2| 243559 + tpg|BK006939.2| 244018 - INS 
 tpg|BK006948.2| 186433 + tpg|BK006948.2| 186037 - INS 
 tpg|BK006939.2| 538867 + tpg|BK006939.2| 538563 - INS 
 tpg|BK006948.2| 202109 + tpg|BK006948.2| 201632 - INS 
 tpg|BK006939.2| 44258 + tpg|BK006939.2| 43704 - INS 
 tpg|BK006948.2| 1069862 + tpg|BK006948.2| 1069899 - INS 
 tpg|BK006948.2| 349582 + tpg|BK006948.2| 349045 - INS 
 tpg|BK006939.2| 45664 + tpg|BK006939.2| 45882 - INS 
 tpg|BK006939.2| 403811 + tpg|BK006939.2| 403045 - INS 
 tpg|BK006948.2| 10773 + tpg|BK006948.2| 10149 - INS 
 tpg|BK006939.2| 366948 + tpg|BK006939.2| 366519 - INS 
 tpg|BK006948.2| 670623 + tpg|BK006948.2| 669921 - INS 
 tpg|BK006939.2| 121690 + tpg|BK006939.2| 121145 - INS 
 tpg|BK006948.2| 366505 + tpg|BK006948.2| 367192 - INS 
 tpg|BK006948.2| 116961 + tpg|BK006948.2| 116811 - INS 
 tpg|BK006939.2| 327177 + tpg|BK006939.2| 326845 - INS 
 tpg|BK006948.2| 428720 + tpg|BK006948.2| 429056 - INS 
 tpg|BK006939.2| 557670 + tpg|BK006939.2| 557663 - INS 
 tpg|BK006948.2| 437268 + tpg|BK006948.2| 436976 - INS 
 tpg|BK006948.2| 15159 + tpg|BK006948.2| 14689 - INS 
 tpg|BK006939.2| 466767 + tpg|BK006939.2| 466913 - INS 
 tpg|BK006939.2| 467961 + tpg|BK006939.2| 467434 - INS 
 tpg|BK006948.2| 772013 + tpg|BK006948.2| 771524 - INS 
 tpg|BK006939.2| 303009 + tpg|BK006939.2| 303629 - INS 
 tpg|BK006948.2| 1008434 + tpg|BK006948.2| 1007703 - INS 
 tpg|BK006939.2| 290881 + tpg|BK006939.2| 291118 - INS 
 tpg|BK006939.2| 24479 + tpg|BK006939.2| 24816 - INS 
 tpg|BK006948.2| 463038 + tpg|BK006948.2| 463712 - INS 
 tpg|BK006939.2| 487237 + tpg|BK006939.2| 486935 - INS 
 tpg|BK006939.2| 23218 + tpg|BK006939.2| 23520 - INS 
 tpg|BK006948.2| 236663 + tpg|BK006948.2| 236519 - INS 
 tpg|BK006948.2| 696632 + tpg|BK006948.2| 696476 - INS 
 tpg|BK006948.2| 958086 + tpg|BK006948.2| 957507 - INS 
 tpg|BK006939.2| 172063 + tpg|BK006939.2| 172379 - INS 
 tpg|BK006948.2| 828335 + tpg|BK006948.2| 828719 - INS 
 tpg|BK006939.2| 213735 + tpg|BK006939.2| 213350 - INS 
 tpg|BK006939.2| 225415 + tpg|BK006939.2| 226041 - INS 
 tpg|BK006948.2| 340396 + tpg|BK006948.2| 339914 - INS 
 tpg|BK006939.2| 289295 + tpg|BK006939.2| 289375 - INS 
 tpg|BK006948.2| 1023922 + tpg|BK006948.2| 1023515 - INS 
 tpg|BK006939.2| 487847 + tpg|BK006939.2| 488199 - INS 
 tpg|BK006939.2| 406464 + tpg|BK006939.2| 407168 - INS 
 tpg|BK006948.2| 1063542 + tpg|BK006948.2| 1063974 - INS 
 tpg|BK006939.2| 11224 + tpg|BK006939.2| 11134 - INS 
 tpg|BK006948.2| 73987 + tpg|BK006948.2| 73767 - INS 
 tpg|BK006939.2| 195411 + tpg|BK006939.2| 195202 - INS 
 tpg|BK006948.2| 966380 + tpg|BK006948.2| 966572 - INS 
 tpg|BK006939.2| 393498 + tpg|BK006939.2| 392772 - INS 
 tpg|BK006939.2| 568581 + tpg|BK006939.2| 568146 - INS 
 tpg|BK006948.2| 262781 + tpg|BK006948.2| 262491 - INS 
 tpg|BK006939.2| 114145 + tpg|BK006939.2| 113931 - INS 
 tpg|BK006948.2| 604088 + tpg|BK006948.2| 603820 - INS 
 tpg|BK006939.2| 520176 + tpg|BK006939.2| 520024 - INS 
 tpg|BK006948.2| 994857 + tpg|BK006948.2| 995020 - INS 
 tpg|BK006939.2| 346987 + tpg|BK006939.2| 346743 - INS 
 tpg|BK006939.2| 134607 + tpg|BK006939.2| 134794 - INS 
 tpg|BK006948.2| 879920 + tpg|BK006948.2| 879445 - INS 
 tpg|BK006939.2| 499370 + tpg|BK006939.2| 499663 - INS 
 tpg|BK006948.2| 574401 + tpg|BK006948.2| 574519 - INS 
 tpg|BK006939.2| 138756 + tpg|BK006939.2| 138976 - INS 
 tpg|BK006939.2| 491285 + tpg|BK006939.2| 491533 - INS 
 tpg|BK006948.2| 1076718 + tpg|BK006948.2| 1076096 - INS 
 tpg|BK006939.2| 299827 + tpg|BK006939.2| 299470 - INS 
 tpg|BK006948.2| 580642 + tpg|BK006948.2| 580417 - INS 
 tpg|BK006939.2| 294258 + tpg|BK006939.2| 294423 - INS 
 tpg|BK006948.2| 89501 + tpg|BK006948.2| 89862 - INS 
 tpg|BK006948.2| 922941 + tpg|BK006948.2| 923221 - INS 
 tpg|BK006948.2| 178509 + tpg|BK006948.2| 177916 - INS 
 tpg|BK006939.2| 272393 + tpg|BK006939.2| 272380 - INS 
 tpg|BK006948.2| 538424 + tpg|BK006948.2| 537790 - INS 
 tpg|BK006939.2| 394277 + tpg|BK006939.2| 394247 - INS 
 tpg|BK006948.2| 648432 + tpg|BK006948.2| 648141 - INS 
 tpg|BK006939.2| 408982 + tpg|BK006939.2| 409725 - INS 
 tpg|BK006948.2| 679665 + tpg|BK006948.2| 680308 - INS 
 tpg|BK006948.2| 39896 + tpg|BK006948.2| 39992 - INS 
 tpg|BK006939.2| 82151 + tpg|BK006939.2| 81580 - INS 
 tpg|BK006939.2| 106134 + tpg|BK006939.2| 106848 - INS 
 tpg|BK006939.2| 93972 + tpg|BK006939.2| 94523 - INS 
 tpg|BK006948.2| 815488 + tpg|BK006948.2| 815599 - INS 
 tpg|BK006939.2| 248756 + tpg|BK006939.2| 248267 - INS 
 tpg|BK006948.2| 931385 + tpg|BK006948.2| 930986 - INS 
 tpg|BK006939.2| 190877 + tpg|BK006939.2| 190535 - INS 
 tpg|BK006948.2| 560769 + tpg|BK006948.2| 560793 - INS 
 tpg|BK006939.2| 87622 + tpg|BK006939.2| 87142 - INS 
 tpg|BK006948.2| 303970 + tpg|BK006948.2| 303364 - INS 
 tpg|BK006948.2| 614704 + tpg|BK006948.2| 614692 - INS 
 tpg|BK006939.2| 438185 + tpg|BK006939.2| 438025 - INS 
 tpg|BK006939.2| 282302 + tpg|BK006939.2| 282927 - INS 
 tpg|BK006948.2| 621914 + tpg|BK006948.2| 621564 - INS 
 tpg|BK006939.2| 28596 + tpg|BK006939.2| 28133 - INS 
 tpg|BK006948.2| 503898 + tpg|BK006948.2| 504125 - INS 
 tpg|BK006948.2| 657435 + tpg|BK006948.2| 657923 - INS 
 tpg|BK006939.2| 151395 + tpg|BK006939.2| 151108 - INS 
 tpg|BK006948.2| 951997 + tpg|BK006948.2| 952622 - INS 
 tpg|BK006939.2| 263163 + tpg|BK006939.2| 262962 - INS 
 tpg|BK006948.2| 1046052 + tpg|BK006948.2| 1045889 - INS 
 tpg|BK006939.2| 140362 + tpg|BK006939.2| 140470 - INS 
 tpg|BK006948.2| 211007 + tpg|BK006948.2| 210375 - INS 
 tpg|BK006939.2| 89786 + tpg|BK006939.2| 89061 - INS 
 tpg|BK006948.2| 859479 + tpg|BK006948.2| 859018 - INS 
 tpg|BK006939.2| 250381 + tpg|BK006939.2| 250472 - INS 
 tpg|BK006939.2| 566303 + tpg|BK006939.2| 566660 - INS 
 tpg|BK006939.2| 476468 + tpg|BK006939.2| 476454 - INS 
 tpg|BK006948.2| 324486 + tpg|BK006948.2| 325190 - INS 
 tpg|BK006948.2| 167374 + tpg|BK006948.2| 167945 - INS 
 tpg|BK006939.2| 537418 + tpg|BK006939.2| 537534 - INS 
 tpg|BK006939.2| 414928 + tpg|BK006939.2| 414269 - INS 
 tpg|BK006948.2| 563824 + tpg|BK006948.2| 563448 - INS 
 tpg|BK006939.2| 179610 + tpg|BK006939.2| 179130 - INS 
 tpg|BK006948.2| 586419 + tpg|BK006948.2| 586104 - INS 
 tpg|BK006939.2| 178860 + tpg|BK006939.2| 178396 - INS 
 tpg|BK006939.2| 39979 + tpg|BK006939.2| 40659 - INS 
 tpg|BK006939.2| 176877 + tpg|BK006939.2| 177508 - INS 
 tpg|BK006939.2| 110329 + tpg|BK006939.2| 110483 - INS 
 tpg|BK006948.2| 405716 + tpg|BK006948.2| 405426 - INS 
 tpg|BK006948.2| 419185 + tpg|BK006948.2| 419148 - INS 
 tpg|BK006939.2| 219222 + tpg|BK006939.2| 219227 - INS 
 tpg|BK006948.2| 221874 + tpg|BK006948.2| 221802 - INS 
 tpg|BK006948.2| 942104 + tpg|BK006948.2| 942357 - INS 
 tpg|BK006939.2| 381406 + tpg|BK006939.2| 381725 - INS 
 tpg|BK006939.2| 379720 + tpg|BK006939.2| 379471 - INS 
 tpg|BK006948.2| 723812 + tpg|BK006948.2| 723471 - INS 
 tpg|BK006939.2| 166412 + tpg|BK006939.2| 166205 - INS 
 tpg|BK006948.2| 946767 + tpg|BK006948.2| 946740 - INS 
 tpg|BK006948.2| 446514 + tpg|BK006948.2| 446262 - INS 
 tpg|BK006948.2| 237225 + tpg|BK006948.2| 237540 - INS 
 tpg|BK006948.2| 714810 + tpg|BK006948.2| 714599 - INS 
 tpg|BK006939.2| 459859 + tpg|BK006939.2| 460359 - INS 
 tpg|BK006939.2| 124294 + tpg|BK006939.2| 124713 - INS 
 tpg|BK006948.2| 84869 + tpg|BK006948.2| 85376 - INS 
 tpg|BK006948.2| 476213 + tpg|BK006948.2| 475784 - INS 
 tpg|BK006939.2| 60951 + tpg|BK006939.2| 60612 - INS 
 tpg|BK006939.2| 315535 + tpg|BK006939.2| 315044 - INS 
 tpg|BK006948.2| 19517 + tpg|BK006948.2| 19691 - INS 
 tpg|BK006939.2| 314790 + tpg|BK006939.2| 314722 - INS 
 tpg|BK006939.2| 132212 + tpg|BK006939.2| 132381 - INS 
 tpg|BK006948.2| 820570 + tpg|BK006948.2| 820366 - INS 
 tpg|BK006948.2| 194784 + tpg|BK006948.2| 194451 - INS 
 tpg|BK006939.2| 297665 + tpg|BK006939.2| 297296 - INS 
 tpg|BK006948.2| 508477 + tpg|BK006948.2| 508812 - INS 
 tpg|BK006939.2| 268121 + tpg|BK006939.2| 267908 - INS 
 tpg|BK006948.2| 108144 + tpg|BK006948.2| 107391 - INS 
 tpg|BK006948.2| 639732 + tpg|BK006948.2| 639476 - INS 
 tpg|BK006939.2| 311414 + tpg|BK006939.2| 311333 - INS 
 tpg|BK006948.2| 1019669 + tpg|BK006948.2| 1020079 - INS 
 tpg|BK006948.2| 605528 + tpg|BK006948.2| 605216 - INS GC
 tpg|BK006948.2| 539488 + tpg|BK006948.2| 539482 - INS 
 tpg|BK006939.2| 68784 + tpg|BK006939.2| 68559 - INS 
 tpg|BK006948.2| 988855 + tpg|BK006948.2| 988630 - INS 
 tpg|BK006939.2| 289916 + tpg|BK006939.2| 290524 - INS 
 tpg|BK006948.2| 587439 + tpg|BK006948.2| 587208 - INS 
 tpg|BK006939.2| 71318 + tpg|BK006939.2| 71534 - INS 
 tpg|BK006939.2| 146991 + tpg|BK006939.2| 147191 - INS 
 tpg|BK006948.2| 282789 + tpg|BK006948.2| 282497 - INS 
 tpg|BK006939.2| 273586 + tpg|BK006939.2| 273273 - INS 
 ref|NC_001224| 20453 + ref|NC_001224| 20238 - INS 
 tpg|BK006948.2| 996654 + tpg|BK006948.2| 996875 - INS 
 tpg|BK006939.2| 257358 + tpg|BK006939.2| 257891 - INS 
 tpg|BK006948.2| 157136 + tpg|BK006948.2| 157659 - INS 
 tpg|BK006939.2| 163259 + tpg|BK006939.2| 163050 - INS 
 tpg|BK006939.2| 86841 + tpg|BK006939.2| 86313 - INS 
 tpg|BK006948.2| 266073 + tpg|BK006948.2| 265520 - INS 
 tpg|BK006939.2| 181855 + tpg|BK006939.2| 181975 - INS 
 tpg|BK006948.2| 851915 + tpg|BK006948.2| 851780 - INS 
 tpg|BK006939.2| 370379 + tpg|BK006939.2| 370380 - INS 
 tpg|BK006948.2| 644579 + tpg|BK006948.2| 644484 - INS 
 tpg|BK006948.2| 831696 + tpg|BK006948.2| 831198 - INS 
 tpg|BK006948.2| 328863 + tpg|BK006948.2| 328296 - INS 
 tpg|BK006939.2| 149246 + tpg|BK006939.2| 149196 - INS 
 tpg|BK006948.2| 499958 + tpg|BK006948.2| 499342 - INS 
 tpg|BK006939.2| 387671 + tpg|BK006939.2| 387683 - INS 
 tpg|BK006948.2| 666839 + tpg|BK006948.2| 667136 - INS 
 tpg|BK006948.2| 802902 + tpg|BK006948.2| 802209 - INS 
 tpg|BK006939.2| 347745 + tpg|BK006939.2| 347455 - INS 
 tpg|BK006948.2| 962148 + tpg|BK006948.2| 962061 - INS 
 tpg|BK006939.2| 265830 + tpg|BK006939.2| 266405 - INS 
 tpg|BK006948.2| 1009019 + tpg|BK006948.2| 1008898 - INS 
 tpg|BK006939.2| 298140 + tpg|BK006939.2| 298492 - INS 
 tpg|BK006948.2| 1057052 + tpg|BK006948.2| 1057162 - INS 
 tpg|BK006939.2| 76789 + tpg|BK006939.2| 76747 - INS 
 tpg|BK006948.2| 785488 + tpg|BK006948.2| 785983 - INS 
 tpg|BK006939.2| 256466 + tpg|BK006939.2| 255893 - INS 
 tpg|BK006948.2| 1052562 + tpg|BK006948.2| 1052740 - INS 
 tpg|BK006948.2| 514408 + tpg|BK006948.2| 513914 - INS 
 tpg|BK006939.2| 454815 + tpg|BK006939.2| 454115 - INS 
 tpg|BK006948.2| 822758 + tpg|BK006948.2| 822841 - INS 
 tpg|BK006939.2| 127852 + tpg|BK006939.2| 127646 - INS 
 tpg|BK006948.2| 35039 + tpg|BK006948.2| 34698 - INS 
 tpg|BK006939.2| 440446 + tpg|BK006939.2| 440128 - INS 
 tpg|BK006948.2| 665695 + tpg|BK006948.2| 665458 - INS 
 tpg|BK006939.2| 173487 + tpg|BK006939.2| 172991 - INS 
 tpg|BK006948.2| 784060 + tpg|BK006948.2| 783448 - INS 
 tpg|BK006939.2| 556513 + tpg|BK006939.2| 555867 - INS 
 tpg|BK006948.2| 114523 + tpg|BK006948.2| 113817 - INS 
 tpg|BK006939.2| 211499 + tpg|BK006939.2| 211109 - INS 
 tpg|BK006948.2| 203861 + tpg|BK006948.2| 203708 - INS 
 tpg|BK006939.2| 398656 + tpg|BK006939.2| 398685 - INS 
 tpg|BK006948.2| 33260 + tpg|BK006948.2| 32926 - INS 
 tpg|BK006939.2| 185365 + tpg|BK006939.2| 185472 - INS 
 tpg|BK006948.2| 472161 + tpg|BK006948.2| 471572 - INS 
 tpg|BK006939.2| 112564 + tpg|BK006939.2| 113191 - INS 
 tpg|BK006948.2| 16735 + tpg|BK006948.2| 16547 - INS 
 tpg|BK006939.2| 175830 + tpg|BK006939.2| 175698 - INS 
 tpg|BK006948.2| 411768 + tpg|BK006948.2| 412229 - INS 
 tpg|BK006939.2| 360702 + tpg|BK006939.2| 360198 - INS 
 tpg|BK006948.2| 406234 + tpg|BK006948.2| 406164 - INS 
 tpg|BK006939.2| 435460 + tpg|BK006939.2| 435071 - INS 
 tpg|BK006939.2| 559264 + tpg|BK006939.2| 558839 - INS 
 tpg|BK006948.2| 17817 + tpg|BK006948.2| 17356 - INS 
 tpg|BK006939.2| 252953 + tpg|BK006939.2| 253603 - INS 
 tpg|BK006948.2| 923562 + tpg|BK006948.2| 923786 - INS 
 tpg|BK006948.2| 239114 + tpg|BK006948.2| 238796 - INS 
 tpg|BK006948.2| 140413 + tpg|BK006948.2| 141154 - INS 
 tpg|BK006948.2| 358576 + tpg|BK006948.2| 358322 - INS 
 tpg|BK006939.2| 255193 + tpg|BK006939.2| 255163 - INS 
 tpg|BK006939.2| 464858 + tpg|BK006939.2| 464950 - INS 
 tpg|BK006948.2| 71518 + tpg|BK006948.2| 70924 - INS 
 tpg|BK006939.2| 142616 + tpg|BK006939.2| 142454 - INS 
 tpg|BK006948.2| 320390 + tpg|BK006948.2| 319973 - INS 
 tpg|BK006939.2| 385283 + tpg|BK006939.2| 385240 - INS 
 tpg|BK006939.2| 228833 + tpg|BK006939.2| 228570 - INS 
 tpg|BK006948.2| 567236 + tpg|BK006948.2| 567467 - INS 
 tpg|BK006939.2| 367845 + tpg|BK006939.2| 367276 - INS 
 tpg|BK006939.2| 390240 + tpg|BK006939.2| 390085 - INS 
 tpg|BK006939.2| 227466 + tpg|BK006939.2| 227051 - INS 
 tpg|BK006948.2| 607011 + tpg|BK006948.2| 606756 - INS 
 tpg|BK006939.2| 130611 + tpg|BK006939.2| 131200 - INS 
 tpg|BK006948.2| 913165 + tpg|BK006948.2| 912599 - INS 
 tpg|BK006948.2| 257161 + tpg|BK006948.2| 256650 - INS 
 tpg|BK006939.2| 323223 + tpg|BK006939.2| 323478 - INS 
 tpg|BK006939.2| 463987 + tpg|BK006939.2| 463653 - INS 
 tpg|BK006948.2| 526224 + tpg|BK006948.2| 525571 - INS 
 tpg|BK006939.2| 304984 + tpg|BK006939.2| 304800 - INS 
 tpg|BK006948.2| 61281 + tpg|BK006948.2| 61333 - INS 
 tpg|BK006939.2| 284602 + tpg|BK006939.2| 285253 - INS 
 tpg|BK006948.2| 645544 + tpg|BK006948.2| 645529 - INS 
 tpg|BK006948.2| 886592 + tpg|BK006948.2| 886023 - INS 
 tpg|BK006939.2| 107724 + tpg|BK006939.2| 107569 - INS 
 tpg|BK006939.2| 292858 + tpg|BK006939.2| 292751 - INS 
 tpg|BK006939.2| 294675 + tpg|BK006939.2| 295433 - INS 
 tpg|BK006939.2| 296348 + tpg|BK006939.2| 296536 - INS 
 tpg|BK006948.2| 207245 + tpg|BK006948.2| 207215 - INS 
 tpg|BK006948.2| 695902 + tpg|BK006948.2| 695221 - INS 
 tpg|BK006939.2| 468699 + tpg|BK006939.2| 468756 - INS 
 tpg|BK006939.2| 306264 + tpg|BK006939.2| 305813 - INS 
 tpg|BK006948.2| 592329 + tpg|BK006948.2| 592084 - INS 
 tpg|BK006939.2| 310150 + tpg|BK006939.2| 309768 - INS 
 tpg|BK006948.2| 529770 + tpg|BK006948.2| 529517 - INS 
 tpg|BK006948.2| 620263 + tpg|BK006948.2| 620865 - INS 
 tpg|BK006939.2| 518132 + tpg|BK006939.2| 517987 - INS 
 tpg|BK006939.2| 338596 + tpg|BK006939.2| 338248 - INS 
 tpg|BK006948.2| 623564 + tpg|BK006948.2| 623242 - INS 
 tpg|BK006939.2| 122162 + tpg|BK006939.2| 122247 - INS 
 tpg|BK006948.2| 746456 + tpg|BK006948.2| 746900 - INS 
 tpg|BK006939.2| 88116 + tpg|BK006939.2| 87919 - INS 
 tpg|BK006948.2| 51679 + tpg|BK006948.2| 51025 - INS 
 tpg|BK006939.2| 544107 + tpg|BK006939.2| 544126 - INS 
 tpg|BK006948.2| 554446 + tpg|BK006948.2| 554315 - INS 
 tpg|BK006948.2| 989471 + tpg|BK006948.2| 989268 - INS 
 tpg|BK006948.2| 775659 + tpg|BK006948.2| 776165 - INS 
 tpg|BK006948.2| 83286 + tpg|BK006948.2| 83033 - INS 
 tpg|BK006948.2| 755611 + tpg|BK006948.2| 755323 - INS 
 tpg|BK006948.2| 135764 + tpg|BK006948.2| 135278 - INS 
 tpg|BK006948.2| 235170 + tpg|BK006948.2| 234786 - INS 
 tpg|BK006948.2| 947713 + tpg|BK006948.2| 947842 - INS 
 tpg|BK006948.2| 779827 + tpg|BK006948.2| 779272 - INS 
 tpg|BK006939.2| 364503 + tpg|BK006939.2| 364602 - INS 
 tpg|BK006939.2| 512230 + tpg|BK006939.2| 511983 - INS 
 tpg|BK006948.2| 474481 + tpg|BK006948.2| 474425 - INS 
 tpg|BK006939.2| 531978 + tpg|BK006939.2| 531707 - INS 
 tpg|BK006948.2| 804693 + tpg|BK006948.2| 804962 - INS 
 tpg|BK006948.2| 340968 + tpg|BK006948.2| 340863 - INS 
 tpg|BK006939.2| 38359 + tpg|BK006939.2| 37948 - INS 
 tpg|BK006948.2| 496705 + tpg|BK006948.2| 496473 - INS 
 tpg|BK006939.2| 408251 + tpg|BK006939.2| 408377 - INS 
 tpg|BK006939.2| 105507 + tpg|BK006939.2| 104960 - INS 
 tpg|BK006948.2| 908275 + tpg|BK006948.2| 908826 - INS 
 tpg|BK006948.2| 857345 + tpg|BK006948.2| 857367 - INS 
 tpg|BK006948.2| 77680 + tpg|BK006948.2| 77802 - INS 
 tpg|BK006939.2| 341788 + tpg|BK006939.2| 342109 - INS 
 tpg|BK006939.2| 276344 + tpg|BK006939.2| 276159 - INS 
 tpg|BK006948.2| 266905 + tpg|BK006948.2| 266792 - INS 
 tpg|BK006939.2| 74651 + tpg|BK006939.2| 74669 - INS 
 tpg|BK006948.2| 99155 + tpg|BK006948.2| 98392 - INS 
 tpg|BK006939.2| 397694 + tpg|BK006939.2| 397443 - INS 
 tpg|BK006939.2| 423280 + tpg|BK006939.2| 422683 - INS 
 tpg|BK006948.2| 385970 + tpg|BK006948.2| 385869 - INS 
 tpg|BK006939.2| 166995 + tpg|BK006939.2| 167120 - INS 
 tpg|BK006939.2| 193474 + tpg|BK006939.2| 192995 - INS 
 tpg|BK006948.2| 452749 + tpg|BK006948.2| 452021 - INS 
 tpg|BK006939.2| 93460 + tpg|BK006939.2| 93264 - INS 
 tpg|BK006948.2| 56291 + tpg|BK006948.2| 55586 - INS 
 tpg|BK006939.2| 138133 + tpg|BK006939.2| 137550 - INS 
 tpg|BK006948.2| 432943 + tpg|BK006948.2| 432912 - INS 
 tpg|BK006939.2| 16036 + tpg|BK006939.2| 15849 - INS 
 tpg|BK006939.2| 384371 + tpg|BK006939.2| 383729 - INS 
 tpg|BK006939.2| 20989 + tpg|BK006939.2| 21694 - INS 
 tpg|BK006948.2| 322913 + tpg|BK006948.2| 322822 - INS 
 tpg|BK006948.2| 766663 + tpg|BK006948.2| 766780 - INS 
 tpg|BK006939.2| 345379 + tpg|BK006939.2| 345955 - INS 
 tpg|BK006939.2| 216797 + tpg|BK006939.2| 217008 - INS 
 tpg|BK006948.2| 388264 + tpg|BK006948.2| 387946 - INS 
 tpg|BK006939.2| 341066 + tpg|BK006939.2| 340978 - INS 
 tpg|BK006939.2| 396621 + tpg|BK006939.2| 396448 - INS 
 tpg|BK006939.2| 514608 + tpg|BK006939.2| 514769 - INS 
 tpg|BK006948.2| 795229 + tpg|BK006948.2| 794480 - INS 
 tpg|BK006948.2| 438490 + tpg|BK006948.2| 437938 - INS 
 tpg|BK006939.2| 506778 + tpg|BK006939.2| 506453 - INS 
 tpg|BK006939.2| 322886 + tpg|BK006939.2| 322325 - INS 
 tpg|BK006948.2| 730582 + tpg|BK006948.2| 730945 - INS 
 tpg|BK006939.2| 56429 + tpg|BK006939.2| 56994 - INS 
 tpg|BK006948.2| 399958 + tpg|BK006948.2| 400306 - INS 
 tpg|BK006939.2| 55099 + tpg|BK006939.2| 55059 - INS 
 tpg|BK006948.2| 935228 + tpg|BK006948.2| 934700 - INS 
 tpg|BK006939.2| 261983 + tpg|BK006939.2| 261598 - INS 
 tpg|BK006939.2| 363054 + tpg|BK006939.2| 363821 - INS 
 tpg|BK006948.2| 753223 + tpg|BK006948.2| 753209 - INS 
 tpg|BK006939.2| 18306 + tpg|BK006939.2| 18690 - INS 
 tpg|BK006948.2| 407962 + tpg|BK006948.2| 408312 - INS 
 tpg|BK006948.2| 411027 + tpg|BK006948.2| 410638 - INS 
 tpg|BK006948.2| 1012782 + tpg|BK006948.2| 1013132 - INS 
 tpg|BK006939.2| 502799 + tpg|BK006939.2| 502778 - INS 
 tpg|BK006939.2| 318719 + tpg|BK006939.2| 318637 - INS 
 tpg|BK006939.2| 246104 + tpg|BK006939.2| 245701 - INS 
 tpg|BK006939.2| 413378 + tpg|BK006939.2| 413229 - INS 
 tpg|BK006948.2| 231921 + tpg|BK006948.2| 231457 - INS 
 tpg|BK006939.2| 351464 + tpg|BK006939.2| 351507 - INS 
 tpg|BK006939.2| 392010 + tpg|BK006939.2| 391750 - INS 
 tpg|BK006939.2| 472394 + tpg|BK006939.2| 472092 - INS 
 tpg|BK006948.2| 728789 + tpg|BK006948.2| 728351 - INS 
 tpg|BK006939.2| 551389 + tpg|BK006939.2| 551779 - INS 
 tpg|BK006948.2| 729789 + tpg|BK006948.2| 729347 - INS 
 tpg|BK006939.2| 153112 + tpg|BK006939.2| 152819 - INS 
 tpg|BK006948.2| 745772 + tpg|BK006948.2| 745992 - INS 
 tpg|BK006939.2| 451651 + tpg|BK006939.2| 451550 - INS 
 tpg|BK006948.2| 968488 + tpg|BK006948.2| 967842 - INS 
 tpg|BK006948.2| 1051605 + tpg|BK006948.2| 1051311 - INS 
 tpg|BK006948.2| 875651 + tpg|BK006948.2| 875169 - INS 
 tpg|BK006948.2| 356411 + tpg|BK006948.2| 356535 - INS 
 tpg|BK006948.2| 889463 + tpg|BK006948.2| 890173 - INS 
 tpg|BK006948.2| 58490 + tpg|BK006948.2| 58229 - INS 
 tpg|BK006948.2| 1054008 + tpg|BK006948.2| 1053718 - INS 
 tpg|BK006948.2| 875986 + tpg|BK006948.2| 876089 - INS 
 tpg|BK006939.2| 548002 + tpg|BK006939.2| 547746 - INS 
 tpg|BK006939.2| 429862 + tpg|BK006939.2| 429697 - INS 
 tpg|BK006939.2| 428681 + tpg|BK006939.2| 427977 - INS 
 tpg|BK006939.2| 421828 + tpg|BK006939.2| 421196 - INS 
 tpg|BK006939.2| 96519 + tpg|BK006939.2| 96575 - INS 
 tpg|BK006948.2| 869969 + tpg|BK006948.2| 869784 - INS 
 tpg|BK006939.2| 419504 + tpg|BK006939.2| 419561 - INS 
 tpg|BK006939.2| 246613 + tpg|BK006939.2| 246302 - INS 
 tpg|BK006948.2| 102201 + tpg|BK006948.2| 101637 - INS 
 tpg|BK006939.2| 111858 + tpg|BK006939.2| 111588 - INS 
 tpg|BK006948.2| 986176 + tpg|BK006948.2| 986202 - INS 
 tpg|BK006939.2| 238921 + tpg|BK006939.2| 238579 - INS 
 tpg|BK006939.2| 95401 + tpg|BK006939.2| 95521 - INS 
 tpg|BK006939.2| 249276 + tpg|BK006939.2| 249030 - INS 
 tpg|BK006948.2| 615580 + tpg|BK006948.2| 615675 - INS 
 tpg|BK006939.2| 475927 + tpg|BK006939.2| 475394 - INS 
 tpg|BK006939.2| 527636 + tpg|BK006939.2| 527613 - INS 
 tpg|BK006948.2| 188051 + tpg|BK006948.2| 187505 - INS 
 tpg|BK006939.2| 521733 + tpg|BK006939.2| 522016 - INS 
 tpg|BK006939.2| 165062 + tpg|BK006939.2| 164670 - INS 
 tpg|BK006948.2| 124605 + tpg|BK006948.2| 125058 - INS 
 tpg|BK006939.2| 357898 + tpg|BK006939.2| 357365 - INS 
 tpg|BK006939.2| 188708 + tpg|BK006939.2| 188160 - INS 
 tpg|BK006939.2| 531178 + tpg|BK006939.2| 530917 - INS 
 tpg|BK006939.2| 186280 + tpg|BK006939.2| 186218 - INS 
 tpg|BK006948.2| 79936 + tpg|BK006948.2| 79690 - INS 
 tpg|BK006939.2| 203645 + tpg|BK006939.2| 203321 - INS 
 tpg|BK006939.2| 533761 + tpg|BK006939.2| 533571 - INS 
 tpg|BK006939.2| 46867 + tpg|BK006939.2| 46838 - INS 
 tpg|BK006948.2| 519289 + tpg|BK006948.2| 519168 - INS 
 tpg|BK006948.2| 277016 + tpg|BK006948.2| 276984 - INS 
 tpg|BK006939.2| 319647 + tpg|BK006939.2| 319623 - INS 
 tpg|BK006939.2| 65994 + tpg|BK006939.2| 65631 - INS 
 tpg|BK006939.2| 10320 + tpg|BK006939.2| 10227 - INS 
 tpg|BK006939.2| 565143 + tpg|BK006939.2| 565010 - INS 
 tpg|BK006939.2| 85391 + tpg|BK006939.2| 85353 - INS 
 tpg|BK006948.2| 650961 + tpg|BK006948.2| 650699 - INS 
 tpg|BK006939.2| 19505 + tpg|BK006939.2| 19270 - INS 
 tpg|BK006948.2| 211932 + tpg|BK006948.2| 212348 - INS 
 tpg|BK006939.2| 425459 + tpg|BK006939.2| 425173 - INS CATATGTTGT
 tpg|BK006948.2| 1047272 + tpg|BK006948.2| 1046882 - INS 
 tpg|BK006939.2| 536644 + tpg|BK006939.2| 537182 - INS 
 tpg|BK006939.2| 216101 + tpg|BK006939.2| 215689 - INS 
 tpg|BK006948.2| 979316 + tpg|BK006948.2| 979198 - INS 
 tpg|BK006939.2| 404305 + tpg|BK006939.2| 404498 - INS 
 tpg|BK006939.2| 77761 + tpg|BK006939.2| 77381 - INS 
 tpg|BK006948.2| 980257 + tpg|BK006948.2| 979689 - INS 
 tpg|BK006948.2| 287099 + tpg|BK006948.2| 287053 - INS 
 tpg|BK006939.2| 148310 + tpg|BK006939.2| 148090 - INS 
 tpg|BK006939.2| 6528 + tpg|BK006939.2| 6646 - INS 
 tpg|BK006948.2| 505830 + tpg|BK006948.2| 505437 - INS 
 tpg|BK006939.2| 169436 + tpg|BK006939.2| 169265 - INS 
 tpg|BK006948.2| 489239 + tpg|BK006948.2| 488962 - INS 
 tpg|BK006939.2| 232534 + tpg|BK006939.2| 232079 - INS 
 tpg|BK006948.2| 661163 + tpg|BK006948.2| 660426 - INS 
 tpg|BK006939.2| 455476 + tpg|BK006939.2| 454980 - INS 
 tpg|BK006939.2| 29608 + tpg|BK006939.2| 29372 - INS 
 tpg|BK006948.2| 62328 + tpg|BK006948.2| 62299 - INS 
 tpg|BK006939.2| 128617 + tpg|BK006939.2| 128664 - INS 
 tpg|BK006939.2| 429210 + tpg|BK006939.2| 428478 - INS 
 tpg|BK006948.2| 664823 + tpg|BK006948.2| 664120 - INS 
 tpg|BK006939.2| 44658 + tpg|BK006939.2| 44499 - INS 
 tpg|BK006948.2| 1010509 + tpg|BK006948.2| 1010720 - INS 
 tpg|BK006939.2| 517181 + tpg|BK006939.2| 516594 - INS 
 tpg|BK006948.2| 467985 + tpg|BK006948.2| 467840 - INS 
 tpg|BK006948.2| 812560 + tpg|BK006948.2| 813175 - INS 
 tpg|BK006939.2| 12446 + tpg|BK006939.2| 13121 - INS 
 tpg|BK006939.2| 286760 + tpg|BK006939.2| 287193 - INS 
 tpg|BK006939.2| 224929 + tpg|BK006939.2| 224178 - INS 
 tpg|BK006939.2| 208443 + tpg|BK006939.2| 207860 - INS 
 tpg|BK006939.2| 233289 + tpg|BK006939.2| 233436 - INS 
 tpg|BK006948.2| 960793 + tpg|BK006948.2| 960751 - INS 
 tpg|BK006939.2| 200630 + tpg|BK006939.2| 200435 - INS 
 tpg|BK006948.2| 310279 + tpg|BK006948.2| 310109 - INS 
 tpg|BK006939.2| 423559 + tpg|BK006939.2| 423333 - INS 
 tpg|BK006939.2| 354351 + tpg|BK006939.2| 355032 - INS 
 tpg|BK006948.2| 484954 + tpg|BK006948.2| 484303 - INS 
 tpg|BK006939.2| 22740 + tpg|BK006939.2| 22227 - INS 
 tpg|BK006939.2| 536065 + tpg|BK006939.2| 535471 - INS 
 tpg|BK006948.2| 484192 + tpg|BK006948.2| 483837 - INS 
 tpg|BK006939.2| 100206 + tpg|BK006939.2| 100736 - INS 
 tpg|BK006948.2| 1015350 + tpg|BK006948.2| 1015122 - INS 
 tpg|BK006939.2| 436006 + tpg|BK006939.2| 436549 - INS 
 tpg|BK006939.2| 306912 + tpg|BK006939.2| 306483 - INS 
 tpg|BK006939.2| 380890 + tpg|BK006939.2| 380160 - INS 
 tpg|BK006948.2| 435445 + tpg|BK006948.2| 435664 - INS 
 tpg|BK006939.2| 184535 + tpg|BK006939.2| 184312 - INS 
 tpg|BK006939.2| 524022 + tpg|BK006939.2| 523783 - INS 
 tpg|BK006939.2| 511687 + tpg|BK006939.2| 511149 - INS 
 tpg|BK006948.2| 770580 + tpg|BK006948.2| 771063 - INS 
 tpg|BK006939.2| 417385 + tpg|BK006939.2| 417566 - INS 
 tpg|BK006939.2| 9524 + tpg|BK006939.2| 9200 - INS 
 tpg|BK006948.2| 824960 + tpg|BK006948.2| 825103 - INS 
 tpg|BK006948.2| 71975 + tpg|BK006948.2| 72522 - INS 
 tpg|BK006948.2| 996068 + tpg|BK006948.2| 995675 - INS 
 tpg|BK006939.2| 530 + tpg|BK006939.2| 321 - INS 
 tpg|BK006939.2| 439293 + tpg|BK006939.2| 439699 - INS 
 ref|NC_001224| 18339 + ref|NC_001224| 18630 - INS 
 tpg|BK006939.2| 135679 + tpg|BK006939.2| 136339 - INS 
 tpg|BK006939.2| 64744 + tpg|BK006939.2| 64778 - INS 
 tpg|BK006948.2| 507240 + tpg|BK006948.2| 506616 - INS 
 tpg|BK006939.2| 443433 + tpg|BK006939.2| 442928 - INS 
 tpg|BK006948.2| 511079 + tpg|BK006948.2| 511827 - INS 
 tpg|BK006948.2| 811275 + tpg|BK006948.2| 811803 - INS 
 tpg|BK006948.2| 323889 + tpg|BK006948.2| 324109 - INS 
 tpg|BK006948.2| 254558 + tpg|BK006948.2| 254567 - INS 
 tpg|BK006948.2| 842934 + tpg|BK006948.2| 842272 - INS 
 tpg|BK006948.2| 855946 + tpg|BK006948.2| 855514 - INS 
 tpg|BK006948.2| 139697 + tpg|BK006948.2| 139386 - INS 
 tpg|BK006948.2| 1000754 + tpg|BK006948.2| 1000982 - INS 
 tpg|BK006948.2| 594415 + tpg|BK006948.2| 594512 - INS 
 tpg|BK006948.2| 999609 + tpg|BK006948.2| 999173 - INS 
 tpg|BK006948.2| 451679 + tpg|BK006948.2| 451398 - INS 
 tpg|BK006948.2| 784696 + tpg|BK006948.2| 784399 - INS 
 tpg|BK006948.2| 593566 + tpg|BK006948.2| 593393 - INS 
 tpg|BK006948.2| 188619 + tpg|BK006948.2| 189256 - INS 
 tpg|BK006948.2| 936316 + tpg|BK006948.2| 936791 - INS 
 tpg|BK006948.2| 752431 + tpg|BK006948.2| 751846 - INS 
 tpg|BK006948.2| 765973 + tpg|BK006948.2| 765616 - INS 
 tpg|BK006948.2| 540946 + tpg|BK006948.2| 541055 - INS 
 tpg|BK006948.2| 84321 + tpg|BK006948.2| 84005 - INS 
 tpg|BK006948.2| 233394 + tpg|BK006948.2| 232899 - INS 
 tpg|BK006948.2| 93776 + tpg|BK006948.2| 93540 - INS 
 tpg|BK006948.2| 790752 + tpg|BK006948.2| 791275 - INS 
 tpg|BK006948.2| 242815 + tpg|BK006948.2| 243065 - INS 
 tpg|BK006948.2| 53958 + tpg|BK006948.2| 53512 - INS 
 tpg|BK006948.2| 672353 + tpg|BK006948.2| 671754 - INS 
 tpg|BK006948.2| 1059831 + tpg|BK006948.2| 1060092 - INS 
 tpg|BK006948.2| 261684 + tpg|BK006948.2| 261156 - INS 
 tpg|BK006948.2| 799902 + tpg|BK006948.2| 799377 - INS 
 tpg|BK006948.2| 86934 + tpg|BK006948.2| 86820 - INS 
 tpg|BK006948.2| 905542 + tpg|BK006948.2| 905122 - INS 
 tpg|BK006948.2| 368994 + tpg|BK006948.2| 368713 - INS 
 tpg|BK006948.2| 983591 + tpg|BK006948.2| 983204 - INS 
 tpg|BK006948.2| 1017544 + tpg|BK006948.2| 1017759 - INS 
 tpg|BK006948.2| 602089 + tpg|BK006948.2| 601831 - INS 
 tpg|BK006948.2| 1407 + tpg|BK006948.2| 1177 - INS 
 tpg|BK006948.2| 699665 + tpg|BK006948.2| 700422 - INS 
 tpg|BK006948.2| 326018 + tpg|BK006948.2| 325748 - INS 
 tpg|BK006948.2| 568330 + tpg|BK006948.2| 568274 - INS 
 tpg|BK006948.2| 569154 + tpg|BK006948.2| 569032 - INS 
 tpg|BK006948.2| 76514 + tpg|BK006948.2| 76443 - INS 
 tpg|BK006948.2| 398518 + tpg|BK006948.2| 398259 - INS 
 tpg|BK006948.2| 18780 + tpg|BK006948.2| 18683 - INS 
 tpg|BK006948.2| 259065 + tpg|BK006948.2| 258790 - INS 
 tpg|BK006948.2| 1003882 + tpg|BK006948.2| 1003739 - INS 
 tpg|BK006948.2| 663980 + tpg|BK006948.2| 663404 - INS 
 tpg|BK006948.2| 683865 + tpg|BK006948.2| 683596 - INS 
 tpg|BK006948.2| 740750 + tpg|BK006948.2| 741322 - INS 
 tpg|BK006948.2| 956468 + tpg|BK006948.2| 956739 - INS 
 tpg|BK006948.2| 824311 + tpg|BK006948.2| 823856 - INS 
 tpg|BK006948.2| 616506 + tpg|BK006948.2| 617008 - INS 
 tpg|BK006948.2| 808480 + tpg|BK006948.2| 807874 - INS 
 tpg|BK006948.2| 763915 + tpg|BK006948.2| 763632 - INS 
 tpg|BK006948.2| 66594 + tpg|BK006948.2| 66809 - INS 
 tpg|BK006948.2| 816772 + tpg|BK006948.2| 816678 - INS 
 tpg|BK006948.2| 1014116 + tpg|BK006948.2| 1014023 - INS 
 tpg|BK006948.2| 749669 + tpg|BK006948.2| 749132 - INS 
 tpg|BK006948.2| 49807 + tpg|BK006948.2| 50029 - INS 
 tpg|BK006948.2| 5314 + tpg|BK006948.2| 5916 - INS 
 tpg|BK006948.2| 850208 + tpg|BK006948.2| 849748 - INS 
 tpg|BK006948.2| 439653 + tpg|BK006948.2| 439064 - INS 
 tpg|BK006948.2| 458188 + tpg|BK006948.2| 457693 - INS 
 tpg|BK006948.2| 674186 + tpg|BK006948.2| 674686 - INS 
 tpg|BK006948.2| 353217 + tpg|BK006948.2| 353100 - INS 
 tpg|BK006948.2| 887395 + tpg|BK006948.2| 887819 - INS 
 tpg|BK006948.2| 507754 + tpg|BK006948.2| 507067 - INS 
 tpg|BK006948.2| 777839 + tpg|BK006948.2| 777721 - INS 
 tpg|BK006948.2| 883936 + tpg|BK006948.2| 884123 - INS 
 tpg|BK006948.2| 880539 + tpg|BK006948.2| 880495 - INS 
 tpg|BK006948.2| 68609 + tpg|BK006948.2| 68961 - INS 
 tpg|BK006948.2| 950643 + tpg|BK006948.2| 949961 - INS 
 tpg|BK006948.2| 633588 + tpg|BK006948.2| 633445 - INS 
 tpg|BK006948.2| 1005346 + tpg|BK006948.2| 1005635 - INS 
 tpg|BK006948.2| 1024469 + tpg|BK006948.2| 1024712 - INS 
 tpg|BK006948.2| 976674 + tpg|BK006948.2| 976163 - INS 
 tpg|BK006948.2| 393900 + tpg|BK006948.2| 393325 - INS 
 tpg|BK006948.2| 99658 + tpg|BK006948.2| 99325 - INS 
 tpg|BK006948.2| 780230 + tpg|BK006948.2| 780138 - INS 
 tpg|BK006948.2| 15724 + tpg|BK006948.2| 15778 - INS 
 tpg|BK006948.2| 179498 + tpg|BK006948.2| 179972 - INS 
 tpg|BK006948.2| 137275 + tpg|BK006948.2| 136914 - INS 
 tpg|BK006948.2| 485843 + tpg|BK006948.2| 486324 - INS 
 tpg|BK006948.2| 150035 + tpg|BK006948.2| 149557 - INS 
 tpg|BK006948.2| 309322 + tpg|BK006948.2| 309652 - INS 
 tpg|BK006948.2| 54861 + tpg|BK006948.2| 54542 - INS 
 tpg|BK006948.2| 832560 + tpg|BK006948.2| 832291 - INS 
 tpg|BK006948.2| 134304 + tpg|BK006948.2| 134220 - INS 
 tpg|BK006948.2| 330543 + tpg|BK006948.2| 330064 - INS 
 tpg|BK006948.2| 555211 + tpg|BK006948.2| 555115 - INS 
 tpg|BK006948.2| 624126 + tpg|BK006948.2| 623785 - INS 
 tpg|BK006948.2| 739331 + tpg|BK006948.2| 739309 - INS 
 tpg|BK006948.2| 160774 + tpg|BK006948.2| 160713 - INS 
 tpg|BK006948.2| 618886 + tpg|BK006948.2| 618639 - INS 
 tpg|BK006948.2| 113441 + tpg|BK006948.2| 112727 - INS 
 tpg|BK006948.2| 581327 + tpg|BK006948.2| 581814 - INS 
 tpg|BK006948.2| 520110 + tpg|BK006948.2| 519667 - INS 
 tpg|BK006948.2| 865086 + tpg|BK006948.2| 864678 - INS 
 tpg|BK006948.2| 978654 + tpg|BK006948.2| 978535 - INS 
 tpg|BK006948.2| 485426 + tpg|BK006948.2| 484896 - INS 
 tpg|BK006948.2| 288206 + tpg|BK006948.2| 287803 - INS 
 tpg|BK006948.2| 154053 + tpg|BK006948.2| 154343 - INS 
 tpg|BK006948.2| 520587 + tpg|BK006948.2| 521021 - INS 
 tpg|BK006948.2| 854411 + tpg|BK006948.2| 854076 - INS 
 tpg|BK006948.2| 958815 + tpg|BK006948.2| 958366 - INS 
 tpg|BK006948.2| 246906 + tpg|BK006948.2| 247060 - INS 
 tpg|BK006948.2| 629870 + tpg|BK006948.2| 629388 - INS 
 tpg|BK006948.2| 60022 + tpg|BK006948.2| 59383 - INS 
 tpg|BK006948.2| 399166 + tpg|BK006948.2| 398986 - INS 
 tpg|BK006948.2| 46946 + tpg|BK006948.2| 47142 - INS 
 tpg|BK006948.2| 500857 + tpg|BK006948.2| 500339 - INS 
 tpg|BK006948.2| 881749 + tpg|BK006948.2| 882456 - INS 
 tpg|BK006948.2| 1024791 + tpg|BK006948.2| 1025423 - INS 
 tpg|BK006948.2| 350051 + tpg|BK006948.2| 349737 - INS 
 tpg|BK006948.2| 220062 + tpg|BK006948.2| 220554 - INS 
 tpg|BK006948.2| 860023 + tpg|BK006948.2| 860073 - INS 
 tpg|BK006948.2| 955944 + tpg|BK006948.2| 955629 - INS 
 tpg|BK006948.2| 91842 + tpg|BK006948.2| 92237 - INS 
 tpg|BK006948.2| 770150 + tpg|BK006948.2| 769892 - INS 
 tpg|BK006948.2| 569753 + tpg|BK006948.2| 570091 - INS 
 tpg|BK006948.2| 23826 + tpg|BK006948.2| 23185 - INS 
 tpg|BK006948.2| 1071493 + tpg|BK006948.2| 1071312 - INS 
 tpg|BK006948.2| 703069 + tpg|BK006948.2| 702858 - INS 
 tpg|BK006948.2| 298398 + tpg|BK006948.2| 297937 - INS 
 tpg|BK006948.2| 935707 + tpg|BK006948.2| 935763 - INS 
 tpg|BK006948.2| 295300 + tpg|BK006948.2| 295256 - INS CA
 tpg|BK006948.2| 268995 + tpg|BK006948.2| 269255 - INS 
 tpg|BK006948.2| 82254 + tpg|BK006948.2| 81578 - INS 
 tpg|BK006948.2| 123948 + tpg|BK006948.2| 123785 - INS 
 tpg|BK006948.2| 345235 + tpg|BK006948.2| 344528 - INS 
 tpg|BK006948.2| 698297 + tpg|BK006948.2| 697586 - INS 
 tpg|BK006948.2| 810556 + tpg|BK006948.2| 810483 - INS 
 tpg|BK006948.2| 252169 + tpg|BK006948.2| 251884 - INS 
 tpg|BK006948.2| 354968 + tpg|BK006948.2| 354260 - INS 
 tpg|BK006948.2| 863897 + tpg|BK006948.2| 864281 - INS 
 tpg|BK006948.2| 109724 + tpg|BK006948.2| 109315 - INS 
 tpg|BK006948.2| 981561 + tpg|BK006948.2| 981204 - INS 
 ref|NC_001224| 61497 + ref|NC_001224| 60929 - INS 
 tpg|BK006948.2| 963870 + tpg|BK006948.2| 964459 - INS 
 tpg|BK006948.2| 977804 + tpg|BK006948.2| 977748 - INS 
 tpg|BK006948.2| 331214 + tpg|BK006948.2| 331160 - INS 
 tpg|BK006948.2| 329330 + tpg|BK006948.2| 328995 - INS 
 tpg|BK006948.2| 589731 + tpg|BK006948.2| 589039 - INS 
 tpg|BK006948.2| 563220 + tpg|BK006948.2| 562856 - INS 
 tpg|BK006948.2| 407152 + tpg|BK006948.2| 406988 - INS 
 tpg|BK006948.2| 902481 + tpg|BK006948.2| 901988 - INS 
 tpg|BK006948.2| 630243 + tpg|BK006948.2| 630032 - INS 
 tpg|BK006948.2| 420661 + tpg|BK006948.2| 420152 - INS 
 tpg|BK006948.2| 941159 + tpg|BK006948.2| 941112 - INS 
 tpg|BK006948.2| 914341 + tpg|BK006948.2| 914825 - INS 
 tpg|BK006948.2| 911609 + tpg|BK006948.2| 911807 - INS 
 tpg|BK006948.2| 728462 + tpg|BK006948.2| 727803 - INS 
 tpg|BK006948.2| 1065778 + tpg|BK006948.2| 1065655 - INS 
 tpg|BK006948.2| 492800 + tpg|BK006948.2| 492599 - INS 
 tpg|BK006948.2| 800562 + tpg|BK006948.2| 800811 - INS 
 tpg|BK006948.2| 476890 + tpg|BK006948.2| 476315 - INS 
 tpg|BK006948.2| 350612 + tpg|BK006948.2| 350642 - INS 
 tpg|BK006948.2| 678369 + tpg|BK006948.2| 678129 - INS 
 tpg|BK006948.2| 190619 + tpg|BK006948.2| 189955 - INS 
 tpg|BK006948.2| 832154 + tpg|BK006948.2| 831650 - INS 
 tpg|BK006948.2| 335821 + tpg|BK006948.2| 335810 - INS 
 tpg|BK006948.2| 183227 + tpg|BK006948.2| 183906 - INS 
 tpg|BK006948.2| 727480 + tpg|BK006948.2| 727309 - INS 
 tpg|BK006948.2| 533016 + tpg|BK006948.2| 533184 - INS 
 tpg|BK006948.2| 951035 + tpg|BK006948.2| 950834 - INS 
 tpg|BK006948.2| 781408 + tpg|BK006948.2| 780661 - INS 
 tpg|BK006948.2| 1078293 + tpg|BK006948.2| 1077952 - INS 
 tpg|BK006948.2| 223160 + tpg|BK006948.2| 222695 - INS 
 tpg|BK006948.2| 336763 + tpg|BK006948.2| 336147 - INS 
 tpg|BK006948.2| 993136 + tpg|BK006948.2| 993160 - INS 
 tpg|BK006948.2| 761827 + tpg|BK006948.2| 761729 - INS 
 tpg|BK006948.2| 686524 + tpg|BK006948.2| 686457 - INS 
 tpg|BK006948.2| 26207 + tpg|BK006948.2| 25830 - INS 
 tpg|BK006948.2| 913891 + tpg|BK006948.2| 913413 - INS 
 tpg|BK006948.2| 20813 + tpg|BK006948.2| 20524 - INS 
 tpg|BK006948.2| 963306 + tpg|BK006948.2| 963701 - INS 
 tpg|BK006948.2| 355616 + tpg|BK006948.2| 354905 - INS 
 tpg|BK006948.2| 37418 + tpg|BK006948.2| 37954 - INS 
 tpg|BK006948.2| 308615 + tpg|BK006948.2| 308340 - INS 
 tpg|BK006948.2| 970137 + tpg|BK006948.2| 969975 - INS 
 tpg|BK006948.2| 625455 + tpg|BK006948.2| 625949 - INS 
 tpg|BK006948.2| 466906 + tpg|BK006948.2| 466796 - INS 
 tpg|BK006948.2| 847896 + tpg|BK006948.2| 847655 - INS 
 ref|NC_001224| 15371 + ref|NC_001224| 14620 - INS 
 ref|NC_001224| 21462 + ref|NC_001224| 21099 - INS 
 ref|NC_001224| 41795 + ref|NC_001224| 41889 - INS 
 ref|NC_001224| 22526 + ref|NC_001224| 22306 - INS 
 tpg|BK006943.2| 385473 + tpg|BK006943.2| 385968 - INS 
 tpg|BK006943.2| 244214 + tpg|BK006943.2| 243472 - INS 
 tpg|BK006943.2| 87628 + tpg|BK006943.2| 88151 - INS 
 tpg|BK006943.2| 357488 + tpg|BK006943.2| 356757 - INS 
 ref|NC_001224| 17847 + ref|NC_001224| 17472 - INS 
 tpg|BK006943.2| 205564 + tpg|BK006943.2| 205934 - INS 
 tpg|BK006943.2| 296476 + tpg|BK006943.2| 296171 - INS 
 tpg|BK006943.2| 696180 + tpg|BK006943.2| 695578 - INS 
 ref|NC_001224| 38521 + ref|NC_001224| 38329 - INS 
 tpg|BK006943.2| 45310 + tpg|BK006943.2| 45241 - INS 
 tpg|BK006943.2| 391715 + tpg|BK006943.2| 391884 - INS 
 tpg|BK006943.2| 76620 + tpg|BK006943.2| 76037 - INS 
 tpg|BK006943.2| 497186 + tpg|BK006943.2| 497748 - INS 
 tpg|BK006943.2| 360922 + tpg|BK006943.2| 361552 - INS 
 tpg|BK006943.2| 647560 + tpg|BK006943.2| 646968 - INS 
 tpg|BK006943.2| 717593 + tpg|BK006943.2| 717496 - INS 
 tpg|BK006943.2| 362990 + tpg|BK006943.2| 362781 - INS 
 tpg|BK006943.2| 151432 + tpg|BK006943.2| 150899 - INS 
 tpg|BK006943.2| 648315 + tpg|BK006943.2| 648828 - INS 
 tpg|BK006943.2| 574687 + tpg|BK006943.2| 574434 - INS 
 tpg|BK006943.2| 349545 + tpg|BK006943.2| 349161 - INS 
 tpg|BK006943.2| 232993 + tpg|BK006943.2| 233406 - INS 
 tpg|BK006943.2| 570354 + tpg|BK006943.2| 569663 - INS 
 ref|NC_001224| 62021 + ref|NC_001224| 61474 - INS 
 tpg|BK006943.2| 169647 + tpg|BK006943.2| 169654 - INS 
 tpg|BK006943.2| 316866 + tpg|BK006943.2| 316640 - INS 
 tpg|BK006943.2| 358180 + tpg|BK006943.2| 357568 - INS 
 tpg|BK006943.2| 608984 + tpg|BK006943.2| 609746 - INS 
 tpg|BK006943.2| 657555 + tpg|BK006943.2| 656868 - INS 
 tpg|BK006943.2| 308337 + tpg|BK006943.2| 308565 - INS 
 tpg|BK006943.2| 521489 + tpg|BK006943.2| 522245 - INS 
 tpg|BK006943.2| 260855 + tpg|BK006943.2| 261057 - INS 
 tpg|BK006943.2| 338171 + tpg|BK006943.2| 338278 - INS 
 tpg|BK006943.2| 525792 + tpg|BK006943.2| 525948 - INS 
 tpg|BK006943.2| 419733 + tpg|BK006943.2| 420090 - INS 
 tpg|BK006943.2| 232256 + tpg|BK006943.2| 231727 - INS 
 tpg|BK006943.2| 84274 + tpg|BK006943.2| 84505 - INS 
 tpg|BK006943.2| 325108 + tpg|BK006943.2| 325024 - INS 
 tpg|BK006943.2| 719097 + tpg|BK006943.2| 718592 - INS 
 tpg|BK006943.2| 250942 + tpg|BK006943.2| 250815 - INS 
 tpg|BK006943.2| 375848 + tpg|BK006943.2| 375713 - INS 
 tpg|BK006943.2| 155442 + tpg|BK006943.2| 156042 - INS 
 tpg|BK006943.2| 158791 + tpg|BK006943.2| 158830 - INS 
 tpg|BK006943.2| 293622 + tpg|BK006943.2| 293050 - INS 
 tpg|BK006943.2| 490340 + tpg|BK006943.2| 490777 - INS 
 tpg|BK006943.2| 561818 + tpg|BK006943.2| 562095 - INS 
 tpg|BK006943.2| 586168 + tpg|BK006943.2| 586433 - INS 
 tpg|BK006943.2| 237978 + tpg|BK006943.2| 238155 - INS 
 ref|NC_001224| 25045 + ref|NC_001224| 24599 - INS 
 tpg|BK006943.2| 241784 + tpg|BK006943.2| 241862 - INS 
 tpg|BK006943.2| 640317 + tpg|BK006943.2| 639708 - INS 
 tpg|BK006943.2| 222943 + tpg|BK006943.2| 222672 - INS 
 tpg|BK006943.2| 705598 + tpg|BK006943.2| 705550 - INS 
 tpg|BK006943.2| 578176 + tpg|BK006943.2| 577904 - INS 
 tpg|BK006943.2| 615382 + tpg|BK006943.2| 615348 - INS 
 tpg|BK006943.2| 663397 + tpg|BK006943.2| 662650 - INS 
 tpg|BK006943.2| 189679 + tpg|BK006943.2| 190054 - INS 
 tpg|BK006943.2| 165404 + tpg|BK006943.2| 165654 - INS 
 tpg|BK006943.2| 87094 + tpg|BK006943.2| 86827 - INS 
 tpg|BK006943.2| 457362 + tpg|BK006943.2| 456592 - INS 
 tpg|BK006943.2| 670006 + tpg|BK006943.2| 670470 - INS 
 tpg|BK006943.2| 465684 + tpg|BK006943.2| 465182 - INS 
 tpg|BK006943.2| 91771 + tpg|BK006943.2| 91565 - INS 
 tpg|BK006943.2| 257255 + tpg|BK006943.2| 257339 - INS 
 tpg|BK006943.2| 571661 + tpg|BK006943.2| 571368 - INS 
 tpg|BK006943.2| 572982 + tpg|BK006943.2| 572622 - INS 
 tpg|BK006943.2| 711263 + tpg|BK006943.2| 710831 - INS 
 tpg|BK006943.2| 60332 + tpg|BK006943.2| 60073 - INS 
 tpg|BK006943.2| 328002 + tpg|BK006943.2| 327383 - INS 
 tpg|BK006943.2| 560772 + tpg|BK006943.2| 560113 - INS 
 tpg|BK006943.2| 94043 + tpg|BK006943.2| 94538 - INS 
 tpg|BK006943.2| 179072 + tpg|BK006943.2| 179326 - INS 
 tpg|BK006943.2| 322093 + tpg|BK006943.2| 321738 - INS 
 tpg|BK006943.2| 675769 + tpg|BK006943.2| 675028 - INS 
 tpg|BK006943.2| 690761 + tpg|BK006943.2| 691057 - INS 
 ref|NC_001224| 39394 + ref|NC_001224| 39528 - INS 
 tpg|BK006943.2| 632304 + tpg|BK006943.2| 632172 - INS 
 tpg|BK006943.2| 468050 + tpg|BK006943.2| 468149 - INS 
 tpg|BK006943.2| 684516 + tpg|BK006943.2| 684414 - INS 
 tpg|BK006943.2| 383210 + tpg|BK006943.2| 382987 - INS 
 tpg|BK006943.2| 50718 + tpg|BK006943.2| 50514 - INS 
 tpg|BK006943.2| 323853 + tpg|BK006943.2| 323864 - INS 
 tpg|BK006943.2| 576940 + tpg|BK006943.2| 576244 - INS 
 tpg|BK006943.2| 157578 + tpg|BK006943.2| 157965 - INS 
 tpg|BK006943.2| 160478 + tpg|BK006943.2| 159952 - INS 
 tpg|BK006943.2| 635035 + tpg|BK006943.2| 634674 - INS 
 tpg|BK006943.2| 139231 + tpg|BK006943.2| 139407 - INS 
 tpg|BK006943.2| 184696 + tpg|BK006943.2| 184391 - INS 
 tpg|BK006943.2| 517861 + tpg|BK006943.2| 518006 - INS 
 tpg|BK006943.2| 626383 + tpg|BK006943.2| 626942 - INS 
 tpg|BK006943.2| 118154 + tpg|BK006943.2| 118449 - INS 
 tpg|BK006943.2| 400570 + tpg|BK006943.2| 400166 - INS 
 tpg|BK006943.2| 715556 + tpg|BK006943.2| 715325 - INS 
 ref|NC_001224| 23281 + ref|NC_001224| 23927 - INS 
 tpg|BK006943.2| 604908 + tpg|BK006943.2| 605567 - INS 
 tpg|BK006943.2| 32857 + tpg|BK006943.2| 33379 - INS 
 tpg|BK006943.2| 410068 + tpg|BK006943.2| 409737 - INS 
 tpg|BK006943.2| 98011 + tpg|BK006943.2| 98233 - INS 
 tpg|BK006943.2| 528712 + tpg|BK006943.2| 528527 - INS 
 tpg|BK006943.2| 504151 + tpg|BK006943.2| 504141 - INS 
 tpg|BK006943.2| 399356 + tpg|BK006943.2| 399053 - INS 
 tpg|BK006943.2| 182250 + tpg|BK006943.2| 181593 - INS 
 tpg|BK006943.2| 459251 + tpg|BK006943.2| 459812 - INS 
 tpg|BK006943.2| 197084 + tpg|BK006943.2| 197082 - INS 
 tpg|BK006943.2| 636947 + tpg|BK006943.2| 636999 - INS 
 tpg|BK006943.2| 72257 + tpg|BK006943.2| 72996 - INS 
 tpg|BK006943.2| 469702 + tpg|BK006943.2| 469632 - INS 
 tpg|BK006943.2| 307079 + tpg|BK006943.2| 306368 - INS 
 tpg|BK006943.2| 284062 + tpg|BK006943.2| 284375 - INS 
 tpg|BK006943.2| 340404 + tpg|BK006943.2| 340070 - INS 
 tpg|BK006943.2| 347208 + tpg|BK006943.2| 347414 - INS 
 tpg|BK006943.2| 540337 + tpg|BK006943.2| 540583 - INS 
 tpg|BK006943.2| 149123 + tpg|BK006943.2| 148820 - INS 
 ref|NC_001224| 37524 + ref|NC_001224| 37098 - INS 
 tpg|BK006943.2| 706786 + tpg|BK006943.2| 707011 - INS 
 tpg|BK006943.2| 628559 + tpg|BK006943.2| 628596 - INS 
 tpg|BK006943.2| 188428 + tpg|BK006943.2| 188116 - INS 
 tpg|BK006943.2| 665999 + tpg|BK006943.2| 666501 - INS 
 tpg|BK006943.2| 674276 + tpg|BK006943.2| 674220 - INS 
 tpg|BK006943.2| 355566 + tpg|BK006943.2| 356087 - INS 
 tpg|BK006943.2| 64429 + tpg|BK006943.2| 63753 - INS 
 tpg|BK006943.2| 178257 + tpg|BK006943.2| 178061 - INS 
 tpg|BK006943.2| 620700 + tpg|BK006943.2| 620852 - INS 
 tpg|BK006943.2| 105665 + tpg|BK006943.2| 105617 - INS 
 tpg|BK006943.2| 721600 + tpg|BK006943.2| 721017 - INS 
 tpg|BK006943.2| 713474 + tpg|BK006943.2| 713582 - INS 
 tpg|BK006943.2| 294099 + tpg|BK006943.2| 293741 - INS 
 tpg|BK006943.2| 539168 + tpg|BK006943.2| 538957 - INS 
 tpg|BK006943.2| 285919 + tpg|BK006943.2| 285958 - INS 
 tpg|BK006943.2| 331270 + tpg|BK006943.2| 331604 - INS 
 tpg|BK006943.2| 389706 + tpg|BK006943.2| 389362 - INS 
 tpg|BK006943.2| 290798 + tpg|BK006943.2| 290568 - INS 
 tpg|BK006943.2| 623487 + tpg|BK006943.2| 623385 - INS 
 ref|NC_001224| 59420 + ref|NC_001224| 59883 - INS 
 tpg|BK006943.2| 299791 + tpg|BK006943.2| 299240 - INS 
 tpg|BK006943.2| 291418 + tpg|BK006943.2| 291849 - INS 
 tpg|BK006943.2| 230735 + tpg|BK006943.2| 230387 - INS 
 tpg|BK006943.2| 415562 + tpg|BK006943.2| 415235 - INS 
 tpg|BK006943.2| 319327 + tpg|BK006943.2| 318865 - INS 
 tpg|BK006943.2| 509936 + tpg|BK006943.2| 510140 - INS 
 tpg|BK006943.2| 353484 + tpg|BK006943.2| 353107 - INS 
 tpg|BK006943.2| 352089 + tpg|BK006943.2| 352540 - INS 
 tpg|BK006943.2| 679632 + tpg|BK006943.2| 679069 - INS 
 tpg|BK006943.2| 304537 + tpg|BK006943.2| 304135 - INS 
 tpg|BK006943.2| 314104 + tpg|BK006943.2| 314405 - INS GGTGTGTG
 tpg|BK006943.2| 566314 + tpg|BK006943.2| 567038 - INS 
 tpg|BK006943.2| 423081 + tpg|BK006943.2| 422461 - INS 
 tpg|BK006943.2| 235548 + tpg|BK006943.2| 235662 - INS 
 tpg|BK006943.2| 438579 + tpg|BK006943.2| 438764 - INS 
 tpg|BK006943.2| 57263 + tpg|BK006943.2| 57213 - INS 
 tpg|BK006943.2| 441270 + tpg|BK006943.2| 441968 - INS 
 tpg|BK006943.2| 426211 + tpg|BK006943.2| 425961 - INS 
 ref|NC_001224| 80165 + ref|NC_001224| 79509 - INS 
 tpg|BK006943.2| 650947 + tpg|BK006943.2| 650489 - INS 
 tpg|BK006943.2| 523885 + tpg|BK006943.2| 523892 - INS 
 tpg|BK006943.2| 273456 + tpg|BK006943.2| 272850 - INS 
 tpg|BK006943.2| 143192 + tpg|BK006943.2| 142769 - INS 
 tpg|BK006943.2| 144021 + tpg|BK006943.2| 143428 - INS 
 tpg|BK006943.2| 668924 + tpg|BK006943.2| 669626 - INS 
 tpg|BK006943.2| 650085 + tpg|BK006943.2| 649806 - INS 
 tpg|BK006943.2| 495109 + tpg|BK006943.2| 494585 - INS 
 tpg|BK006943.2| 520173 + tpg|BK006943.2| 520057 - INS 
 tpg|BK006943.2| 234384 + tpg|BK006943.2| 234784 - INS 
 tpg|BK006943.2| 384224 + tpg|BK006943.2| 383984 - INS 
 tpg|BK006943.2| 621684 + tpg|BK006943.2| 621210 - INS 
 tpg|BK006943.2| 373961 + tpg|BK006943.2| 373325 - INS 
 tpg|BK006943.2| 388209 + tpg|BK006943.2| 388980 - INS 
 tpg|BK006943.2| 401185 + tpg|BK006943.2| 401005 - INS 
 tpg|BK006943.2| 600680 + tpg|BK006943.2| 600455 - INS 
 tpg|BK006943.2| 443444 + tpg|BK006943.2| 443163 - INS 
 tpg|BK006943.2| 239025 + tpg|BK006943.2| 239080 - INS 
 tpg|BK006943.2| 601369 + tpg|BK006943.2| 601256 - INS 
 tpg|BK006943.2| 81623 + tpg|BK006943.2| 81555 - INS 
 tpg|BK006943.2| 711836 + tpg|BK006943.2| 712313 - INS 
 tpg|BK006943.2| 38972 + tpg|BK006943.2| 38870 - INS 
 tpg|BK006943.2| 263040 + tpg|BK006943.2| 263025 - INS 
 tpg|BK006943.2| 210201 + tpg|BK006943.2| 209700 - INS 
 tpg|BK006943.2| 363797 + tpg|BK006943.2| 364528 - INS 
 tpg|BK006943.2| 180811 + tpg|BK006943.2| 181101 - INS 
 ref|NC_001224| 74421 + ref|NC_001224| 73751 - INS 
 tpg|BK006943.2| 74038 + tpg|BK006943.2| 73790 - INS 
 tpg|BK006943.2| 395709 + tpg|BK006943.2| 396266 - INS 
 tpg|BK006943.2| 655247 + tpg|BK006943.2| 654835 - INS 
 tpg|BK006943.2| 112648 + tpg|BK006943.2| 112441 - INS 
 tpg|BK006943.2| 224129 + tpg|BK006943.2| 223604 - INS 
 tpg|BK006943.2| 427120 + tpg|BK006943.2| 427699 - INS 
 tpg|BK006943.2| 345074 + tpg|BK006943.2| 344505 - INS 
 tpg|BK006943.2| 564904 + tpg|BK006943.2| 564914 - INS 
 tpg|BK006943.2| 726993 + tpg|BK006943.2| 727095 - INS 
 tpg|BK006943.2| 658581 + tpg|BK006943.2| 658725 - INS 
 tpg|BK006943.2| 336601 + tpg|BK006943.2| 335836 - INS 
 tpg|BK006943.2| 432144 + tpg|BK006943.2| 431739 - INS GTTGTCC
 tpg|BK006943.2| 141112 + tpg|BK006943.2| 141814 - INS 
 ref|NC_001224| 40721 + ref|NC_001224| 41177 - INS 
 tpg|BK006943.2| 556091 + tpg|BK006943.2| 555742 - INS 
 tpg|BK006943.2| 329446 + tpg|BK006943.2| 330201 - INS 
 tpg|BK006943.2| 150005 + tpg|BK006943.2| 150313 - INS 
 tpg|BK006943.2| 245503 + tpg|BK006943.2| 244907 - INS 
 tpg|BK006943.2| 249669 + tpg|BK006943.2| 249744 - INS 
 tpg|BK006943.2| 454237 + tpg|BK006943.2| 454394 - INS 
 tpg|BK006943.2| 254540 + tpg|BK006943.2| 254552 - INS 
 tpg|BK006943.2| 295017 + tpg|BK006943.2| 295253 - INS 
 tpg|BK006943.2| 288031 + tpg|BK006943.2| 287734 - INS 
 tpg|BK006943.2| 672864 + tpg|BK006943.2| 672256 - INS 
 tpg|BK006943.2| 486420 + tpg|BK006943.2| 486353 - INS 
 tpg|BK006943.2| 487382 + tpg|BK006943.2| 487161 - INS 
 tpg|BK006943.2| 54031 + tpg|BK006943.2| 54361 - INS 
 tpg|BK006943.2| 529469 + tpg|BK006943.2| 529691 - INS 
 tpg|BK006943.2| 271193 + tpg|BK006943.2| 271679 - INS 
 tpg|BK006943.2| 221649 + tpg|BK006943.2| 221879 - INS 
 tpg|BK006943.2| 546038 + tpg|BK006943.2| 546734 - INS 
 tpg|BK006943.2| 280558 + tpg|BK006943.2| 280766 - INS 
 tpg|BK006943.2| 501875 + tpg|BK006943.2| 502299 - INS 
 tpg|BK006943.2| 307537 + tpg|BK006943.2| 307035 - INS 
 tpg|BK006943.2| 624224 + tpg|BK006943.2| 623967 - INS 
 ref|NC_001224| 25835 + ref|NC_001224| 25241 - INS 
 tpg|BK006943.2| 378815 + tpg|BK006943.2| 378277 - INS 
 tpg|BK006943.2| 394324 + tpg|BK006943.2| 393762 - INS 
 tpg|BK006943.2| 172964 + tpg|BK006943.2| 172978 - INS 
 tpg|BK006943.2| 493091 + tpg|BK006943.2| 493517 - INS 
 tpg|BK006943.2| 495616 + tpg|BK006943.2| 496157 - INS 
 tpg|BK006943.2| 499286 + tpg|BK006943.2| 499484 - INS 
 tpg|BK006943.2| 511133 + tpg|BK006943.2| 511489 - INS 
 tpg|BK006943.2| 23051 + tpg|BK006943.2| 22569 - INS 
 tpg|BK006943.2| 55859 + tpg|BK006943.2| 55271 - INS 
 tpg|BK006943.2| 545603 + tpg|BK006943.2| 545532 - INS 
 tpg|BK006943.2| 90270 + tpg|BK006943.2| 89965 - INS 
 tpg|BK006943.2| 125740 + tpg|BK006943.2| 126000 - INS 
 tpg|BK006943.2| 403696 + tpg|BK006943.2| 403462 - INS 
 tpg|BK006943.2| 135406 + tpg|BK006943.2| 134847 - INS 
 tpg|BK006943.2| 119689 + tpg|BK006943.2| 119340 - INS 
 tpg|BK006943.2| 208422 + tpg|BK006943.2| 207928 - INS 
 tpg|BK006943.2| 380347 + tpg|BK006943.2| 379903 - INS 
 tpg|BK006943.2| 326560 + tpg|BK006943.2| 326367 - INS 
 tpg|BK006943.2| 432638 + tpg|BK006943.2| 433242 - INS 
 tpg|BK006943.2| 334790 + tpg|BK006943.2| 334553 - INS 
 tpg|BK006943.2| 49505 + tpg|BK006943.2| 49255 - INS 
 tpg|BK006943.2| 404686 + tpg|BK006943.2| 405326 - INS 
 ref|NC_001224| 40307 + ref|NC_001224| 39968 - INS 
 tpg|BK006943.2| 587654 + tpg|BK006943.2| 587793 - INS 
 tpg|BK006943.2| 610761 + tpg|BK006943.2| 611474 - INS 
 tpg|BK006943.2| 78961 + tpg|BK006943.2| 78199 - INS 
 tpg|BK006943.2| 26260 + tpg|BK006943.2| 26366 - INS 
 tpg|BK006943.2| 436331 + tpg|BK006943.2| 436622 - INS 
 tpg|BK006943.2| 444875 + tpg|BK006943.2| 445105 - INS 
 tpg|BK006943.2| 140535 + tpg|BK006943.2| 141094 - INS 
 tpg|BK006943.2| 724781 + tpg|BK006943.2| 724565 - INS 
 tpg|BK006943.2| 643419 + tpg|BK006943.2| 642719 - INS 
 tpg|BK006943.2| 598649 + tpg|BK006943.2| 598301 - INS 
 tpg|BK006943.2| 204969 + tpg|BK006943.2| 204480 - INS 
 tpg|BK006943.2| 585567 + tpg|BK006943.2| 585091 - INS 
 tpg|BK006943.2| 557016 + tpg|BK006943.2| 556928 - INS 
 tpg|BK006943.2| 342176 + tpg|BK006943.2| 342750 - INS 
 tpg|BK006943.2| 514295 + tpg|BK006943.2| 513573 - INS 
 tpg|BK006943.2| 444134 + tpg|BK006943.2| 444583 - INS 
 tpg|BK006943.2| 406884 + tpg|BK006943.2| 406572 - INS 
 tpg|BK006943.2| 573640 + tpg|BK006943.2| 573788 - INS 
 ref|NC_001224| 75622 + ref|NC_001224| 75049 - INS 
 tpg|BK006943.2| 350203 + tpg|BK006943.2| 350020 - INS 
 tpg|BK006943.2| 435556 + tpg|BK006943.2| 435185 - INS 
 tpg|BK006943.2| 455686 + tpg|BK006943.2| 455113 - INS 
 tpg|BK006943.2| 317530 + tpg|BK006943.2| 317253 - INS 
 tpg|BK006943.2| 111350 + tpg|BK006943.2| 111213 - INS 
 tpg|BK006943.2| 32192 + tpg|BK006943.2| 32116 - INS 
 tpg|BK006943.2| 470844 + tpg|BK006943.2| 470472 - INS 
 tpg|BK006943.2| 264016 + tpg|BK006943.2| 263851 - INS 
 tpg|BK006943.2| 270291 + tpg|BK006943.2| 270033 - INS 
 tpg|BK006943.2| 137490 + tpg|BK006943.2| 137125 - INS 
 tpg|BK006943.2| 515153 + tpg|BK006943.2| 515309 - INS 
 tpg|BK006943.2| 524716 + tpg|BK006943.2| 525451 - INS 
 tpg|BK006943.2| 268767 + tpg|BK006943.2| 269274 - INS 
 tpg|BK006943.2| 430703 + tpg|BK006943.2| 430057 - INS 
 tpg|BK006943.2| 430148 + tpg|BK006943.2| 429630 - INS 
 tpg|BK006943.2| 97368 + tpg|BK006943.2| 97075 - INS 
 tpg|BK006943.2| 582274 + tpg|BK006943.2| 582384 - INS 
 tpg|BK006943.2| 211927 + tpg|BK006943.2| 211343 - INS 
 tpg|BK006943.2| 411584 + tpg|BK006943.2| 411272 - INS 
 tpg|BK006943.2| 397209 + tpg|BK006943.2| 396993 - INS 
 tpg|BK006943.2| 406158 + tpg|BK006943.2| 405896 - INS 
 tpg|BK006943.2| 171977 + tpg|BK006943.2| 171591 - INS 
 tpg|BK006943.2| 170800 + tpg|BK006943.2| 170487 - INS 
 tpg|BK006943.2| 370873 + tpg|BK006943.2| 371406 - INS 
 tpg|BK006943.2| 180157 + tpg|BK006943.2| 180576 - INS 
 tpg|BK006943.2| 298302 + tpg|BK006943.2| 298196 - INS 
 tpg|BK006943.2| 44176 + tpg|BK006943.2| 44430 - INS 
 tpg|BK006943.2| 82562 + tpg|BK006943.2| 82844 - INS 
 tpg|BK006943.2| 425495 + tpg|BK006943.2| 425401 - INS 
 tpg|BK006943.2| 315828 + tpg|BK006943.2| 315752 - INS 
 tpg|BK006943.2| 339054 + tpg|BK006943.2| 339102 - INS 
 tpg|BK006943.2| 599086 + tpg|BK006943.2| 599434 - INS 
 tpg|BK006943.2| 579399 + tpg|BK006943.2| 579763 - INS 
 tpg|BK006943.2| 446798 + tpg|BK006943.2| 446652 - INS 
 tpg|BK006943.2| 136319 + tpg|BK006943.2| 136584 - INS 
 tpg|BK006943.2| 452154 + tpg|BK006943.2| 452145 - INS 
 tpg|BK006943.2| 654371 + tpg|BK006943.2| 654113 - INS 
 ref|NC_001224| 28941 + ref|NC_001224| 28759 - INS 
 tpg|BK006943.2| 417432 + tpg|BK006943.2| 417067 - INS 
 tpg|BK006943.2| 164328 + tpg|BK006943.2| 164373 - INS 
 tpg|BK006943.2| 492052 + tpg|BK006943.2| 491611 - INS 
 tpg|BK006943.2| 505873 + tpg|BK006943.2| 505350 - INS 
 tpg|BK006943.2| 277819 + tpg|BK006943.2| 277645 - INS 
 tpg|BK006943.2| 276451 + tpg|BK006943.2| 275704 - INS 
 tpg|BK006943.2| 215830 + tpg|BK006943.2| 215360 - INS 
 tpg|BK006943.2| 258844 + tpg|BK006943.2| 258284 - INS 
 tpg|BK006943.2| 638763 + tpg|BK006943.2| 639206 - INS 
 tpg|BK006943.2| 226229 + tpg|BK006943.2| 225949 - INS 
 tpg|BK006943.2| 95979 + tpg|BK006943.2| 95530 - INS 
 ref|NC_001224| 58864 + ref|NC_001224| 58494 - INS 
 tpg|BK006943.2| 367783 + tpg|BK006943.2| 368457 - INS 
 tpg|BK006943.2| 285177 + tpg|BK006943.2| 284858 - INS 
 tpg|BK006943.2| 332633 + tpg|BK006943.2| 332368 - INS 
 tpg|BK006943.2| 193569 + tpg|BK006943.2| 194040 - INS 
 tpg|BK006943.2| 462079 + tpg|BK006943.2| 461484 - INS 
 tpg|BK006943.2| 255489 + tpg|BK006943.2| 255266 - INS 
 tpg|BK006943.2| 561150 + tpg|BK006943.2| 560805 - INS 
 tpg|BK006943.2| 704587 + tpg|BK006943.2| 704684 - INS 
 tpg|BK006943.2| 583592 + tpg|BK006943.2| 583214 - INS 
 tpg|BK006943.2| 613011 + tpg|BK006943.2| 613138 - INS 
 tpg|BK006943.2| 723190 + tpg|BK006943.2| 722761 - INS 
 tpg|BK006943.2| 209641 + tpg|BK006943.2| 209259 - INS 
 tpg|BK006943.2| 85386 + tpg|BK006943.2| 85436 - INS 
 tpg|BK006943.2| 680866 + tpg|BK006943.2| 680922 - INS 
 tpg|BK006943.2| 703775 + tpg|BK006943.2| 703436 - INS 
 tpg|BK006943.2| 107426 + tpg|BK006943.2| 107182 - INS 
 tpg|BK006943.2| 116251 + tpg|BK006943.2| 116533 - INS 
 tpg|BK006943.2| 671680 + tpg|BK006943.2| 671341 - INS 
 tpg|BK006943.2| 228078 + tpg|BK006943.2| 228129 - INS 
 tpg|BK006943.2| 126884 + tpg|BK006943.2| 126503 - INS 
 tpg|BK006943.2| 147716 + tpg|BK006943.2| 147526 - INS 
 tpg|BK006943.2| 102602 + tpg|BK006943.2| 103038 - INS 
 tpg|BK006943.2| 439585 + tpg|BK006943.2| 439713 - INS 
 tpg|BK006943.2| 162514 + tpg|BK006943.2| 162531 - INS 
 tpg|BK006943.2| 686946 + tpg|BK006943.2| 687305 - INS 
 tpg|BK006943.2| 183429 + tpg|BK006943.2| 183260 - INS 
 ref|NC_001224| 13832 + ref|NC_001224| 14132 - INS 
 tpg|BK006943.2| 596502 + tpg|BK006943.2| 597193 - INS 
 tpg|BK006943.2| 652082 + tpg|BK006943.2| 652315 - INS 
 tpg|BK006943.2| 40660 + tpg|BK006943.2| 40668 - INS 
 tpg|BK006943.2| 516837 + tpg|BK006943.2| 516495 - INS 
 tpg|BK006943.2| 125222 + tpg|BK006943.2| 125111 - INS 
 tpg|BK006943.2| 653203 + tpg|BK006943.2| 653416 - INS 
 tpg|BK006943.2| 595250 + tpg|BK006943.2| 594787 - INS 
 tpg|BK006943.2| 282123 + tpg|BK006943.2| 281669 - INS 
 tpg|BK006943.2| 450404 + tpg|BK006943.2| 450080 - INS 
 tpg|BK006943.2| 176230 + tpg|BK006943.2| 175682 - INS 
 tpg|BK006943.2| 374433 + tpg|BK006943.2| 373931 - INS 
 tpg|BK006943.2| 369422 + tpg|BK006943.2| 368949 - INS 
 tpg|BK006943.2| 196279 + tpg|BK006943.2| 196084 - INS 
 tpg|BK006943.2| 68153 + tpg|BK006943.2| 67989 - INS 
 tpg|BK006943.2| 417891 + tpg|BK006943.2| 417745 - INS 
 tpg|BK006943.2| 372513 + tpg|BK006943.2| 372095 - INS 
 tpg|BK006943.2| 630237 + tpg|BK006943.2| 630174 - INS 
 tpg|BK006943.2| 635604 + tpg|BK006943.2| 635350 - INS 
 tpg|BK006943.2| 489725 + tpg|BK006943.2| 490101 - INS 
 tpg|BK006943.2| 682142 + tpg|BK006943.2| 682090 - INS 
 tpg|BK006943.2| 682874 + tpg|BK006943.2| 682974 - INS 
 tpg|BK006943.2| 273896 + tpg|BK006943.2| 274391 - INS 
 tpg|BK006943.2| 562793 + tpg|BK006943.2| 563241 - INS 
 tpg|BK006943.2| 507193 + tpg|BK006943.2| 506777 - INS 
 tpg|BK006943.2| 345625 + tpg|BK006943.2| 345129 - INS 
 tpg|BK006943.2| 680067 + tpg|BK006943.2| 680281 - INS 
 tpg|BK006943.2| 341083 + tpg|BK006943.2| 340710 - INS 
 tpg|BK006943.2| 661689 + tpg|BK006943.2| 661817 - INS 
 ref|NC_001224| 62392 + ref|NC_001224| 61819 - INS 
 tpg|BK006943.2| 668372 + tpg|BK006943.2| 668783 - INS 
 tpg|BK006943.2| 346467 + tpg|BK006943.2| 345897 - INS 
 tpg|BK006943.2| 74970 + tpg|BK006943.2| 74301 - INS 
 tpg|BK006943.2| 195542 + tpg|BK006943.2| 194956 - INS 
 tpg|BK006943.2| 466224 + tpg|BK006943.2| 466710 - INS 
 tpg|BK006943.2| 533241 + tpg|BK006943.2| 533628 - INS 
 tpg|BK006943.2| 492524 + tpg|BK006943.2| 492297 - INS 
 tpg|BK006943.2| 549980 + tpg|BK006943.2| 549495 - INS 
 tpg|BK006943.2| 282663 + tpg|BK006943.2| 282227 - INS 
 tpg|BK006943.2| 602224 + tpg|BK006943.2| 601885 - INS 
 tpg|BK006943.2| 664163 + tpg|BK006943.2| 663726 - INS 
 tpg|BK006943.2| 145697 + tpg|BK006943.2| 145822 - INS 
 tpg|BK006943.2| 35594 + tpg|BK006943.2| 36311 - INS 
 tpg|BK006943.2| 226937 + tpg|BK006943.2| 226525 - INS 
 tpg|BK006943.2| 633393 + tpg|BK006943.2| 633620 - INS 
 tpg|BK006943.2| 591735 + tpg|BK006943.2| 591769 - INS 
 tpg|BK006943.2| 622517 + tpg|BK006943.2| 622229 - INS 
 tpg|BK006943.2| 467357 + tpg|BK006943.2| 467287 - INS 
 tpg|BK006943.2| 115093 + tpg|BK006943.2| 114650 - INS 
 tpg|BK006943.2| 447725 + tpg|BK006943.2| 447504 - INS 
 tpg|BK006943.2| 702638 + tpg|BK006943.2| 702833 - INS 
 tpg|BK006943.2| 697001 + tpg|BK006943.2| 696402 - INS 
 tpg|BK006943.2| 564075 + tpg|BK006943.2| 564203 - INS 
 tpg|BK006943.2| 61777 + tpg|BK006943.2| 61669 - INS 
 tpg|BK006943.2| 256206 + tpg|BK006943.2| 256776 - INS 
 tpg|BK006943.2| 593545 + tpg|BK006943.2| 594094 - INS 
 tpg|BK006943.2| 279802 + tpg|BK006943.2| 280123 - INS 
 tpg|BK006943.2| 220070 + tpg|BK006943.2| 220246 - INS 
 tpg|BK006943.2| 145042 + tpg|BK006943.2| 144505 - INS 
 tpg|BK006943.2| 167254 + tpg|BK006943.2| 166654 - INS 
 tpg|BK006943.2| 319908 + tpg|BK006943.2| 319723 - INS 
 tpg|BK006943.2| 686154 + tpg|BK006943.2| 685633 - INS 
 tpg|BK006943.2| 246525 + tpg|BK006943.2| 246001 - INS 
 tpg|BK006943.2| 424028 + tpg|BK006943.2| 423974 - INS 
 tpg|BK006943.2| 182983 + tpg|BK006943.2| 182527 - INS 
 tpg|BK006943.2| 168547 + tpg|BK006943.2| 168797 - INS 
 tpg|BK006943.2| 595737 + tpg|BK006943.2| 595931 - INS 
 tpg|BK006943.2| 618057 + tpg|BK006943.2| 618026 - INS 
 tpg|BK006943.2| 692725 + tpg|BK006943.2| 692786 - INS 
 tpg|BK006943.2| 351323 + tpg|BK006943.2| 350947 - INS 
 tpg|BK006943.2| 279313 + tpg|BK006943.2| 278680 - INS 
 tpg|BK006943.2| 644202 + tpg|BK006943.2| 643682 - INS 
 tpg|BK006943.2| 309656 + tpg|BK006943.2| 309226 - INS 
 tpg|BK006943.2| 568141 + tpg|BK006943.2| 567852 - INS 
 tpg|BK006943.2| 418703 + tpg|BK006943.2| 418812 - INS 
 tpg|BK006943.2| 124632 + tpg|BK006943.2| 124400 - INS 
 tpg|BK006943.2| 240156 + tpg|BK006943.2| 240635 - INS 
 tpg|BK006943.2| 360118 + tpg|BK006943.2| 359889 - INS 
 tpg|BK006943.2| 51608 + tpg|BK006943.2| 51338 - INS 
 tpg|BK006943.2| 506547 + tpg|BK006943.2| 506329 - INS 
 tpg|BK006943.2| 697401 + tpg|BK006943.2| 698051 - INS 
 tpg|BK006943.2| 457783 + tpg|BK006943.2| 457341 - INS 
 tpg|BK006943.2| 722359 + tpg|BK006943.2| 721731 - INS 
 tpg|BK006943.2| 716124 + tpg|BK006943.2| 716801 - INS 
 tpg|BK006943.2| 602870 + tpg|BK006943.2| 603418 - INS 
 tpg|BK006943.2| 29365 + tpg|BK006943.2| 30092 - INS 
 tpg|BK006943.2| 41591 + tpg|BK006943.2| 41569 - INS 
 tpg|BK006943.2| 604249 + tpg|BK006943.2| 604561 - INS 
 tpg|BK006943.2| 34194 + tpg|BK006943.2| 34674 - INS 
 tpg|BK006943.2| 387553 + tpg|BK006943.2| 387620 - INS 
 tpg|BK006943.2| 507723 + tpg|BK006943.2| 507439 - INS 
 tpg|BK006943.2| 578710 + tpg|BK006943.2| 578838 - INS 
 tpg|BK006943.2| 266333 + tpg|BK006943.2| 266711 - INS 
 tpg|BK006943.2| 311208 + tpg|BK006943.2| 311762 - INS 
 tpg|BK006943.2| 416067 + tpg|BK006943.2| 416089 - INS 
 tpg|BK006943.2| 69861 + tpg|BK006943.2| 69861 - INS 
 tpg|BK006943.2| 225032 + tpg|BK006943.2| 224639 - INS 
 tpg|BK006943.2| 625623 + tpg|BK006943.2| 625939 - INS 
 tpg|BK006943.2| 227327 + tpg|BK006943.2| 227623 - INS 
 tpg|BK006943.2| 79408 + tpg|BK006943.2| 78985 - INS 
 tpg|BK006943.2| 289156 + tpg|BK006943.2| 288795 - INS CAG
 tpg|BK006943.2| 21666 + tpg|BK006943.2| 21555 - INS 
 tpg|BK006943.2| 729284 + tpg|BK006943.2| 728926 - INS 
 tpg|BK006943.2| 541842 + tpg|BK006943.2| 541484 - INS 
 tpg|BK006943.2| 509069 + tpg|BK006943.2| 508533 - INS 
 tpg|BK006943.2| 728411 + tpg|BK006943.2| 727705 - INS 
 tpg|BK006943.2| 173987 + tpg|BK006943.2| 173504 - INS 
 tpg|BK006943.2| 394963 + tpg|BK006943.2| 394434 - INS 
 tpg|BK006943.2| 606443 + tpg|BK006943.2| 606101 - INS 
 tpg|BK006943.2| 174540 + tpg|BK006943.2| 174440 - INS 
 tpg|BK006943.2| 694263 + tpg|BK006943.2| 694173 - INS 
 tpg|BK006943.2| 229000 + tpg|BK006943.2| 229142 - INS 
 tpg|BK006943.2| 471526 + tpg|BK006943.2| 470917 - INS 
 tpg|BK006943.2| 354850 + tpg|BK006943.2| 355275 - INS 
 tpg|BK006943.2| 464296 + tpg|BK006943.2| 464664 - INS 
 tpg|BK006943.2| 232555 + tpg|BK006943.2| 232681 - INS 
 tpg|BK006943.2| 186132 + tpg|BK006943.2| 185749 - INS 
 tpg|BK006943.2| 315192 + tpg|BK006943.2| 314951 - INS 
 tpg|BK006943.2| 547786 + tpg|BK006943.2| 548239 - INS 
 tpg|BK006943.2| 369964 + tpg|BK006943.2| 369888 - INS 
 tpg|BK006943.2| 160952 + tpg|BK006943.2| 160634 - INS 
 tpg|BK006943.2| 631369 + tpg|BK006943.2| 630683 - INS 
 tpg|BK006943.2| 472306 + tpg|BK006943.2| 472127 - INS 
 tpg|BK006943.2| 689933 + tpg|BK006943.2| 690400 - INS 
 tpg|BK006943.2| 199423 + tpg|BK006943.2| 199832 - INS 
 ref|NC_001224| 43807 + ref|NC_001224| 44009 - INS 
 tpg|BK006943.2| 310721 + tpg|BK006943.2| 310472 - INS 
 tpg|BK006943.2| 95435 + tpg|BK006943.2| 95134 - INS 
 tpg|BK006943.2| 414444 + tpg|BK006943.2| 414509 - INS 
 tpg|BK006943.2| 52653 + tpg|BK006943.2| 51956 - INS 
 tpg|BK006943.2| 153541 + tpg|BK006943.2| 153107 - INS 
 tpg|BK006943.2| 185535 + tpg|BK006943.2| 185029 - INS 
 tpg|BK006943.2| 702031 + tpg|BK006943.2| 702062 - INS 
 tpg|BK006943.2| 259311 + tpg|BK006943.2| 259271 - INS 
 tpg|BK006943.2| 512746 + tpg|BK006943.2| 512190 - INS 
 ref|NC_001224| 42704 + ref|NC_001224| 42376 - INS 
 ref|NC_001224| 29640 + ref|NC_001224| 29168 - INS 
 ref|NC_001224| 26396 + ref|NC_001224| 25996 - INS 
 ref|NC_001224| 50711 + ref|NC_001224| 50961 - INS 
 ref|NC_001224| 76245 + ref|NC_001224| 75571 - INS 
 ref|NC_001224| 7926 + ref|NC_001224| 7236 - INS 
 ref|NC_001224| 65886 + ref|NC_001224| 65859 - INS 
 ref|NC_001224| 1172 + ref|NC_001224| 469 - INS 
 ref|NC_001224| 31582 + ref|NC_001224| 30829 - INS 
 ref|NC_001224| 34143 + ref|NC_001224| 34899 - INS 
 ref|NC_001224| 57438 + ref|NC_001224| 57783 - INS 
 ref|NC_001224| 62893 + ref|NC_001224| 62251 - INS 
 ref|NC_001224| 84363 + ref|NC_001224| 84095 - INS 
 ref|NC_001224| 36313 + ref|NC_001224| 36552 - INS 
 ref|NC_001224| 26829 + ref|NC_001224| 26434 - INS 
 ref|NC_001224| 81725 + ref|NC_001224| 81616 - INS 
 ref|NC_001224| 45307 + ref|NC_001224| 44596 - INS TATT
 ref|NC_001224| 35717 + ref|NC_001224| 35762 - INS 
 ref|NC_001224| 2319 + ref|NC_001224| 2186 - INS 
 ref|NC_001224| 33493 + ref|NC_001224| 32922 - INS 
 ref|NC_001224| 27763 + ref|NC_001224| 28303 - INS 
 ref|NC_001224| 80808 + ref|NC_001224| 80406 - INS 
 ref|NC_001224| 54021 + ref|NC_001224| 53735 - INS 
 ref|NC_001224| 5394 + ref|NC_001224| 4964 - INS 
 ref|NC_001224| 63541 + ref|NC_001224| 63461 - INS 
 ref|NC_001224| 77225 + ref|NC_001224| 76609 - INS 
 ref|NC_001224| 47056 + ref|NC_001224| 47803 - INS 
 ref|NC_001224| 46088 + ref|NC_001224| 45493 - INS 
 ref|NC_001224| 72552 + ref|NC_001224| 73220 - INS 
 ref|NC_001224| 64747 + ref|NC_001224| 64496 - INS 
 ref|NC_001224| 53354 + ref|NC_001224| 53156 - INS 
 ref|NC_001224| 78044 + ref|NC_001224| 77527 - INS 
 ref|NC_001224| 3101 + ref|NC_001224| 2698 - INS 
 ref|NC_001224| 67461 + ref|NC_001224| 67224 - INS 
 ref|NC_001224| 68517 + ref|NC_001224| 68404 - INS 
 ref|NC_001224| 56328 + ref|NC_001224| 56679 - INS 
 ref|NC_001224| 84927 + ref|NC_001224| 84647 - INS 
 ref|NC_001224| 12660 + ref|NC_001224| 12316 - INS 
 ref|NC_001224| 6340 + ref|NC_001224| 6184 - INS 
 ref|NC_001224| 46379 + ref|NC_001224| 45865 - INS 
 ref|NC_001224| 55623 + ref|NC_001224| 55042 - INS 
 ref|NC_001224| 69559 + ref|NC_001224| 69749 - INS 
 ref|NC_001224| 50014 + ref|NC_001224| 49774 - INS 
 ref|NC_001224| 83100 + ref|NC_001224| 82673 - INS 
 ref|NC_001224| 85779 + ref|NC_001224| 85528 - INS 
 ref|NC_001224| 9101 + ref|NC_001224| 8759 - INS 
 ref|NC_001224| 56670 + ref|NC_001224| 57141 - INS 
 ref|NC_001224| 70982 + ref|NC_001224| 70592 - INS 
 ref|NC_001224| 3700 + ref|NC_001224| 4017 - INS 
 ref|NC_001224| 8266 + ref|NC_001224| 7839 - INS 
 ref|NC_001224| 71384 + ref|NC_001224| 71279 - INS 
