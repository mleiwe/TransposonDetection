 tpg|BK006937.2| 148614 + tpg|BK006937.2| 148181 - INS CTTCAGTCTTTTTCCATAGGCGAGTCCACAGGGACTACAAAGTTCCCTGTTTTGGTCGGGTCCACTACGCCATTGAATTGTCCAAGTGTCTTTACATTTAGAGCATTCCTTTATCTCACCATTTGGGAGGATTGTTTGTCTCTTTTCTCTTTTAGGACGACTAGTAGTCTTTTTGCTGTATTTCTTCGTAATACTGGCAGACCGACTAGTTCCTTGTGCACAACTATGGTAGCCTTCAAGATTGTTTGCTTCTTGGCTAGTCGTACGTCTCTCGGAATTGCATGCACTAGTTACACGATTCTTTGAGGGTGTAATTTTGTTGGAATAAAAATCAACTATCATCTACTAACTAGTATTTACGTTACTAGTATATTATCATATACGGTGTTAGAAGATGACGCAAATGATGAGAAATAGTCATCTAAATTAGTGGAAGCTGAAACGCAAGGATTGATAATGTAATAGGATCAATGAATATTAACATATAAAACGATGATAATAATATTTATAGAATTGTGTAGAATTGCAGATTCCCTTTTATGGATTCCTAAATCCTTGAGGAGAACTTCTAGTATATTCTGTATACCTAATATTATAGCCTTTATCAACAATGGAATCCCAACAATTATCTCAACATTCACCCATTTCTCATGGTAGCGCCTGTGCTTCGGTTACTTCTAAGGAAGTCCACACAAATCAAGATCCGTTAGACGTTTCAGCTTCCAAAACAGAAGAATGTGAGAAGGCTTCCACTAAGGCTAACTCTCAACAGACAACAACACCTGCTTCATCAGCTGTTCCAGAG
 tpg|BK006935.2| 158649 + tpg|BK006935.2| 158104 - INS GCGCATAGCGAATTTTCTCTCATTTGCATTCAAGTTTGAGTTTGAATGCAGCATATCAGGGACACCAGCATTGCTGGCGTTTGTTTGATTGGCAACATTACCACTGTCAGTTATATCTTCGTCTTTTAAGGTTTCATTTGGATGCTCTGAGAAATAGTTATCCAAAAAAGTACTAGTTTGGTTGACCATATCAGCACGCGACTGGACCAACTCAAAGTCATCTACTAAAAGAACGTATTTCTTTCTTTCCCTGACAATAGCAGGTTCTGCAATTATCACGCGAATGATATCACCCCTTTGTAG
 tpg|BK006935.2| 205910 + tpg|BK006935.2| 205727 - INS CCACAGAAATGACTACTATCACTGGCACCAACGGTGTACCAACTGACGAAACCATCATTGTTGTCAAAACACCAACAACTGCTAGCACCATCATAACTACAACTGAGCCATGGACTGGCACTTTCACCTCTACGTCTACTGAGATGACTACTATCACTGGCACCAACGGTGTACCAACTGACGAAACCATCATTGTTGTCAAAACACCAACAACTGCTAGCACCATCATAACTACGACCGAACCATGGACCGGTACTTTCACATCTACATCCACAGAAATGACTACTGTCACCGGTACCAACGGTCAACCAACTGACGAAACTGTGATTGTTATCAGAACCCCAACTAGTGAAGGTTTGGTTACAACCACCACTGAACCATGGACTGGTACTTTTACCTCTACATCTACTGAGATGACCACCGTCACCGGTACCAACGGTCAACCAACTGACGAAACTGTGATTGTTATCAGAACCCCAACTAGTGAAGGTTTGGTTACAACCACCACTGAACCATGGACTGGTACTTTTACCTCTACATCTACTGAGATGACCACCGTCACCGGTACCAACGGTCAACCAACTGACGAAACTGTGATTGTTATCAGAACCCCAACTAGTGAAGGTTTGGTTACAACCACCACTGAACCATGGACTGGTACTTTTACCTCTACATCTACTGAGATGACCACCATCACTGGAACC
 tpg|BK006935.2| 68008 + tpg|BK006935.2| 67502 - INS ATCTGTATCCTTCAATATGGCCATCGTACAGAAAGCGTATCAAATCAGTGTCTTGAACGAGAGTAAAAGGGAGATGCAATGGAATGTAAGAAATGCTATGGGTCAGAAAAGAAATGCAGAGGAGTTAAACCGAATGAGGAAATGCAATGGATACGTTAAATTGGAGATGTGAGATTGCGACTGGGACTCGGATGGATGCTTGCTTTTGGAGGCTAGTACAGAGAAAAAAGAGGGAGAAAAGAAAAGAGAAATAGAAAAAGGTTGGTTTAAGTCGGCAGAGGAGACTACTCGGGCAATTCGTTTCCTAATGGGCATAGTCCTCTTTCCTCAGAAATCCATTTGACTGGCAGACTCAGTAGT
 tpg|BK006937.2| 59938 + tpg|BK006937.2| 60389 - INS CTTGGACACCGCATGCGTTTCTACACAATGCCGGTAACGATGCCTACTATACCCTGCATTTGTTCATGAAGTTTTGCGATGTTAATTTCAGGAAAATAAGCGGCATGGACGATGTTCTTAAAGTAATGGGCCAAGTAAAAGTTTGGGGAGAACGAGACGTACGAGAGCCTAAAGTGGTGCCCATGTCGTATGCCATCTCCATCG
 tpg|BK006934.2| 502041 + tpg|BK006934.2| 501848 - INS GGTTAGAGAGTAGATGTCCTTATCATATATTATTCCAAGTCGTGGTTACAGGATATCACTAACTTAAGAAAAGTTATTATTTTTTACTTTAGTGTCCTTATCGATCAGTCGCTCTTTCGCCAACTAGCCGCCAATTGCAAAAGCCGATAAGCTTATTTCCCCTCAAGCCGTCAACAAGAACTACAGCAATAACAAAGAGAGTGAATGCAATAAAGGTGTGCGCAACAGTGTAAAATGATACTAAAGCTTGTACACTGTTTAGTTGCTCTTACAGGATTAATCTTTGCAAAGCCGTATCA
 tpg|BK006934.2| 127725 + tpg|BK006934.2| 128105 - INS AAATCAATTGAAAAAGGCAAACGAAAATGGGTTTTCAAGCTGCGTACCGCCAAGCATCACGAAGAAGGAGTTAATAGATGCATGTGGATTTAATCCAAGAGATATGAATAATGAAAGGCAAATTTACGCTCTTCAAGACACCAATTTAGGATTGGTGGCTACCGCGGAGATACCTTTGGCAGGTCTAGGGGCAAACAAAGTTCTAGAGTTAAACTCGGGAGAATGTTCTAAGAAACTAGTTGGAGTAAGTAGATGTTACAGAGCTGAGGCAGGTGCCAGGGGAAAAGATACGAAAGGTCTCTATCG
 tpg|BK006934.2| 562642 + tpg|BK006934.2| 562380 - INS GCTGTAGGGCTAAAGAACAGGATTTCATTTTCATTTTTTTTTTTAATTTCGGTCAGAAAGCCGGGTAAGGAGTGACAGCGAGAGTAAAGATAGATGTGAAAAGTGTGGGTGTGGTGTGTGGGTGTGTGGGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGTGTGTGTGTGGGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGTGGGTGTGTGTGGGTGTGGTGTGTGTGGGTG
 tpg|BK006934.2| 306684 + tpg|BK006934.2| 306317 - INS TTCCAGAAGCTTTAAGTCACTCCTTCATACCGGAATTAGCTAAACAGTTTATCCATTTGTGTTACGACGAAACATATTACAACAAAAGAGGCGGTGTCTTGGGTATAAAAGTTCTCATTGATAATGTTAAGTCGTCCTCAGTTTTCCTAAAAAAGTATCAGTATAACCTAGCCAATGGTCTATTATTTGTGCTGAAGGACACTCAGAGCGAGGCCCCATCTGCTATAACAGATAGCGCTGAGAAATTACTAATAGATCTATTAAGTATTACGTTCGCGGATGTAAAAGA
 tpg|BK006938.2| 1525555 + tpg|BK006938.2| 1525394 - INS GGTGGGATTAGAGTGGTAGAGTAAGTATGTGTGTATTATTTACGATCATTTGTTAGCGTTTCAATAGTGGTGGGTAGAACAATAGTATGGTGAGTAGTAGATGGGAGATGGTAGGGTAAGTGGTAGTGGAGTTGGATATGGGTAATTGGAGGGTAACGGTTATGGTGGACGGTCGGTTGGTGGTAGTACACAGGGAGATGGATGGTGGTTGGGGTGGTATAGTTGAATGAGTCAGGGTAACGAGTGGGGAGGTAGGGTAATGGAGGGTAAGTTGAGAGACAGGTTGGTCAGGGTTGGATTGTGTTAGTGTTAGGGTTAGGGTTGTGTGTGGTGTGGTGTGTGGGTGTGGTGTGTGGTGTGGTGGGTGTGGGTGTGTGGGTGTGGGTGTGTGTGGGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGTGTGGTGTGTGGGTGTGGTGTGGTGTGGTGTGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGTGTGGTGTGTGGGTGTGGTGTGGTGTGGTGTGTGTGGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGTGGTGTGTGTGTGGTGTGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGGGTGTGGTGTGGTGTGTGTGGGTGTGGTGTGGTGTGTATATATATGTCACTGTATTGCATGCTGGATGGTGTTAGACAAGGCCGTAGGGACATATAGCAT
 tpg|BK006941.2| 1063098 + tpg|BK006941.2| 1063583 - INS CTTTTTCTTAATAAATAAGGGAGAAATGTACAGTTAGAATCGTAGAATTATCCACATATCCCTATCTTCAAGATCTGTCGTACTTAAATGCCTCCATAGGTTGCAATCCCCATTTAGCCAACATTGCCTTGTCTTCGTCCCAACCGTTACACATTGTCGTCAGCATTTTCTTACCGGTGAAGATACTGTTACAACCTGCCATGAAACAGACAAATTGCTCTGTTTCTTTCATTGTATAACGACCAGCGGCAAGTCTTATAATGGCCTTTGGCATAACT
 tpg|BK006941.2| 341317 + tpg|BK006941.2| 340565 - INS AAATGATTTAGACAAGTTTTCTTTACCCTATGATGATCCTATTGGAGTTATTTTCCAACTATATGCTGCGAATGAAAATACGGAGAAGCTCTATAAGGAGGTTAGACAAAGAACCAACGCTTTAGATGTTCAGTTTTGCTGGTACTTGATTCAAACATTGAGATTTAATGGAACACGCGTTTTTTCGAAGGAAACTAGCGATGAGGCTACATTCGCATTTGCCGCTCAACTTGAATTTGCACAATTACATGGCCACTCTCTTTTTGTTTCTTGCTTTTTAAATGATGACAAGGCAGCAGAAGATACCATAAAAAGGCTTGTTATGCGTGAAATAACATTGTTAAGAGCCTCTACCAATGATCACATTTTAAAT
 tpg|BK006940.2| 78884 + tpg|BK006940.2| 78878 - INS CTTTTATCGGTAGCCTTAGACTCTAGAAGAGGTAAGATGTGCTTACATTTGTTGCCCAGTTTGTTTAATATCGATACTTCGAATTTGGCGTTATGTGGCGGGATATCGAAATCTAGTGCTAGACATTTAATGGCATATGTATCCGACCTATAAATCCTAGCAGTTCTAGTAGATTTGACCAACTGACAGTGTGTAATGTCTATAC
 tpg|BK006941.2| 62775 + tpg|BK006941.2| 62751 - INS CCCTTCGACTTAGCATTGAAAGAATGGACATCATTAATCAAGTTGTGAAGCTGGTCAATAAAGAGGGTTCTGAGTTTAATCATACTGTGGACTTGAAGAACTATGATAAATTGATTCTAGTGGAATGTTTTAAGAGCAATATCGGAATGTGTGTAGTCGATGGGGATTATAAAACCAAATATCGTAAATACAACGTTCAACAGCTTTATGAATCGAAATTCCGAAAGGATGAAGATAAGAGTGTAAAACAATAATCATATATGAAACAGAATAGATATTTTATATAAGTATATACG
 tpg|BK006938.2| 77718 + tpg|BK006938.2| 77310 - INS TTTTATCAGGATGAATTCCTGCAGGAACAGGCTTGTTGTCTGTTCCAGAGGTTTGAGCTGCAGTGGCGGTAGTTTTGGCGATTTTCTTTTGGTTGCCGTCGTTAATCATCTTTGTCAACCTCTCTTTACGTTCTTCATCCAACTTGATGTTTTTGTTTTTCAATTTTTCTAGACGCTCTTGACTGTTACCACCTCCGCCAACAGTTAGCTCGACATTGATCTTCTTCTCTTTCAGTAAGGTCCCATGTTGTAATAAGGCAATGTCCATACGTCTTTGAATGCCGGTGCGATCTTTGTCAGCATCGAATTCCAAAAATGCAATACCTTTGTCAGCTCTGAGGCGGATCTGGTCGGGTGAACTATTTTTAAAATGGTTTTGCAATTCAACAGCAGTGATGTCTCTAGGTAAGCTACCGACAAAGACAATAAATC
 tpg|BK006941.2| 34872 + tpg|BK006941.2| 34152 - INS CGATATTCAATTGAAGAAAGTGAAAGACACGATGAAACTGCTATTGAAACCCAAGAATTTGATGAAAATGATTGTCTTTCATCTAAGGCGGATATTAATACATCATTAGCTCCTCAAAAGAGATCTTTCATCGATAATGAACTAATGTCCATGTTAGTCACCAAAAAAAAAATAAAGAAGGACAAGGATGTTAGTGACACCGGTATATCTTCCACTTCATACTTGATAAATTCTGGGACATATGCAAATTCTCATATTGAAATTCCTACCTCTAATTC
 tpg|BK006941.2| 265627 + tpg|BK006941.2| 265469 - INS CCAGCAGATGATCTCAATATGTCCCGATAGGCCAATTTTGCCACCAGATAGTTCGATGGCATTTTATTTTTAGTCCTTTTGAAAGCAATATCATAAAATAGATATAGTTCTCCATGATGTTCGGGTCAGTCGCTCCGAAGCGTAACCTAGTATAATAAATAGTTCATTGCAGAAAATAACGAAAGAAATGGTGGAATACGATCTGTTATATCTAAACTAAAGCTAACTAACGGAATAAGCAAATACGAATCGACCGCTAATTTAACAAATATGGTTTTAGCAATGGAAAGTAGAGTGGCACCGGAAATTCCTGGGCTCATTCAACCTGGGAATGTC
 tpg|BK006946.2| 924426 + tpg|BK006946.2| 923710 - INS AGGTAGAAGAACAGTATGGTGAGTAGCAGATGGTGGATGGTAGAGGAATAGCAGGGTAAGTGGTAGTGGAGTTGGATATGGGTAATTGGAGGGTAACGGTTATGGTGCACGATGGGTTGGTGGTAGCAAGTAGAGAGATGGATGGTGGTTGGAGCGGTATGGTTGAAGGGGACAGGGTAACGAGTGGGGAGGTAGCGTAATGGAGGGTAAGTTAAGAGACATGCTAAATCAGGGTAAGAATAGGGTAGGGTTAGGGTAGGGTTAGGGTAGTGTTAGGGTGTGGGTGTGGTGTGTGTGTGTGGGTGTGGTGTGTGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGTGTGGGTGTGTGGGTGTGTGTGTGGGTGTGTGGGTGTGTGGGTGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGGTGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGTGGGTGTGTGTGTGTGGGTGTGTGTGGGTGTGGGTGTGGGTGTGGGTGTGTGGGTGTGGTG
 tpg|BK006938.2| 1120247 + tpg|BK006938.2| 1119801 - INS GCTAAAGCCTGGACAAGCTAAGGAATAATTTGAATTCGCTGATTGAAGAGATCAATGAAAGGTCAGAAACTCAGACAAAAGATGAGAACAACACTGCGAATGACCAATACTCGTCTATTTTGGGGAATTCATTCAATAAATCTTCAAATGACACCATAGAACACGCTGCTGATATAACTGATGGAAATAACACAGAAT
 tpg|BK006946.2| 230739 + tpg|BK006946.2| 230616 - INS CGGCCTTTGCGACCGCCTTTGTCTCTGTCTTGATAGCTGCGCCATTTGTTATGGTCATGAAAGTAGCGCCCGATTTACCTTTCTTATTGGGCGCCTCATTAGTGCTTTTCTTTGTACCAAAGAAGTCTTCGATCGTAGTTTGCTTTCTCTTTCGAGCCACCGTCATAACTGAATTTGTTGGCAATCTTCTCATGCACCACATGTATGTGAACGGCTTGTGTACAGCTTCTGATAATATATATCATTATGGATGAATTACGCGT
 tpg|BK006938.2| 130052 + tpg|BK006938.2| 129519 - INS GTTTCTGTTTCTTACTCCAAATACACTAATGTCTTGAACAAGTTTTATGATTCCAATTACCCTGAATTTCCTGTTTTAAGAGATCGTATGAAGGAAATTCTATCAAACGCTGAAGAATTAGAACAAGTTGTTCAATTAGTTGGTAAATCGGCCTTGTCTGATAGTGATAAGATTACTTTGGATGTTGCCACTTTAATCAAGGAAGATTTCTTGCAACAAAATGGTTACTCCACTTATGATGCTTTCTGTCCAATTTGGAAGACATTTGATATGATGAGAGCCTTCATCTCGTATCATGACGAAGCTCAAAAAGCTGTTGCTAATGGTGCCAACTGGTCAAAACTAGCTGACTCTACTGGTGACGTTAAGCATGCCGTTTCTTCATCTAAATTTTTTGAACCAAGCAGGGGTGAAAAGGAAGTCCATTGCGAATTCGAAAAATTGTTGAGCAC
 tpg|BK006946.2| 601517 + tpg|BK006946.2| 601569 - INS CCTTGTCCAAAGAGAGATTTATGTGAACTGCTTTTGTTTGAAGATAGGTATCAACACCACTTTGCCCCAGTTCTCTACCAATACCACTCATTTTAAACCCGCCAAAAGGAACGGTAACATCTTCATCGTTAGATGAGTTGATCCAAACAGTTCCTGCTTTAATATCGCGAGCAAACATGTGCGCTTTCTTGACATCTTTTGTGAAGACCGCAGAGGCGAGCCCGTAGCAAGTATCATTAGCCAGCTTCAGAGCGTCATCATAATTTGTGAACTTGCTAACAACCACAACCGGGCCAAATATCTCATCCTGTAACAGTTTCGATGTTTGCGGGACATCAGTGAAGATGGTTGGGGGAATGAAGTAGCCTTTAGCTCCACCAATAGGAAATTCAGAGGTCTGGAACATGTCCAACTTTTCCTCCCTTGTACCACGTTCTATGTAACTTTTGATGCGGTCATACTGTGTACTTG
 tpg|BK006946.2| 485787 + tpg|BK006946.2| 485020 - INS TATATGCAGATGGTCCAAGATTACTAAAAGAATTAAGTGACCGTGCTCAAATACCTGTCACCACTACTTTACAAGGTTTAGGTTCATTCGACCAAGAAGATCCAAAATCATTGGATATGCTTGGTATGCACGGTTGTGCTACTGCCAACCTGGCAGTGCAAAATGCCGACTTGATAATTGCAGTTGGTGCTAGATTCGACGACCGTGTCACTGGTAATATTTCTAAATTCGCTCCAGAAGCTCGTCGTGCAGCTGCCGAGGGTAGAGGTGGTATTATTCATTGCGAGGTTAGTCCAAAAAACATAAACAAGGTTGTTCAAACTCAAATAGCAGTGGAAGGTGATGC
 tpg|BK006946.2| 434993 + tpg|BK006946.2| 435501 - INS GGGTTAAATCAGAGGTATTCTCTCATGTGGTGAAGTCCATCAATATCAAGGGTTATTATGTTGGTAACAGAGCTGATACGAGAGAAGCCTTAGACTTCTTTAGCAGAGGTTTGATCAAATCACCAATCAAAATTGTTGGATTATCTGAATTACCAAAGGTTTATGACTTGATGGAAAAGGGCAAGATTTTGGGTAGATACGTCGTCGATACTAGTAAATAATAGCGTGTTACGCACCCAAACTTTTTATGAAAGTCTTTGTTTATAATGATGAGGTTTATAAATATATAGTGGAGCAAAGATTAATCACTAAATCAAGAAGCAGTACCAGTATTTTTTCTATATCAAGTAGTGATAATGGAAATAGCCCAAATTTGGCTTCCGTCGACACAGAGAACGTTTGAGAGACATTATCACCATCAAGCATCGAGC
 tpg|BK006946.2| 5646 + tpg|BK006946.2| 5443 - INS CGTACAAGGTTACTTCCTAGATGCTATATGTCCCTACGGCCTTGTCTAACACCATCCAGCATGCAATACAGTGACATATATATACACACACCACACCCACACACCACACCCACACACACACCACACCCACACACCCACACACCACACCCACACACCCACACCCACACCCACACCCACACACCACACCCACACCCACCCACCACACCC
 tpg|BK006947.3| 23364 + tpg|BK006947.3| 23151 - INS TTTAGAATGGTACCATTCACAACTAATATAGCCTCTGCTGGTTCCTTTAGTAACCTCTTTAGTAACCTCTTTAGTGAAATGGTTCTTGCTGGCTCTATTATTTTCCTAATTCGGACGCGCTGGCTCCGCGCCGTGAGGAAAAACAGCAGGCTGACAAGGGACTAATTTACTGACACTTTCGGCTGACACTTCCGAAAAGGTACTCAAGCTTTTATGAGTAAGATGCTGGTTTGATGCTAAGAATACGATTTAGTACTTCCTTTTTAATGTGGCTTGTTTTTTTTTTATTCGTCCATAAC
 tpg|BK006936.2| 813184 + tpg|BK006936.2| 813033 - INS GTGGTTGGGAGTGGTATGGTTGAATGAGACAGGGTAACGAGTGGGGAGGTAGGGTAATGGAGGGTAGGTTTGGAGACAGGTTCATCAGGGTTAGAATAGGGTACTGTTAGGATTGTGTTAGGGTGTGTGGGTGTGGGTGTGGTGTGTGTGGGTGTGGTGTGTGGGTGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGTGTGTGGGTGTGGGTGTGGGTGTGGGTGTGTGGGTGTGGTGTGTGGTGTGGGTGTGGTGTGTGTGGGTG
 tpg|BK006945.2| 11460 + tpg|BK006945.2| 11207 - INS GTCTAACACCATCCAGCATGCAATACAGTGACATATATATACCACACCCACACACCACACCCACACACACACACCCACACACACACACCACACCCACACACACACACCCACACCACACCCACACACACACCCACACCACACCCACACCCACACACCCACACACACCACACCCACACACCACACCCACACCACACCCACACTCTCTTACATCTACCTCTACTCTCGCTGTCACTCCTTACCCGGCTTTCTGACCGAAATTAAAAAAAATGAAAATGAAACCCTGCTCTTTAGCCCTACAGCACTTCTACAT
 tpg|BK006945.2| 85698 + tpg|BK006945.2| 86151 - INS TGGTCATTGCCCGAGGCCAGATTGTACGCAATGGTCATTGCAGGTACCGTTTTCCCTATTGGTATCTTATGGTTCTGTTGGACGGGCTACTATCCTCACAAGATTCATTGGATGGTCCCCACAGTAGGAGGGGCCTTCATCGGGTTCGGTTTAATGGGTATTTTCTTGCCATGTTTAAACTATATCATTGAATCGTATCTATTGTTGGCAGCTTCTGCCGTCGCAGCAAACACTTTCATGAGGTCTGCATTTGGTGCATGCTTCCCATTGTTTGCAGGATATATGT
 tpg|BK006936.2| 93422 + tpg|BK006936.2| 93571 - INS TTGCTGTCAGAGAAAAAATAGTTTTAAAGGAGACGGTGAACCTTTACCTTCCTTGATATGCAAATATTTTTCAGCTTTTCCTAAAACTAAACATTCTCGACTTTTTTTTAGAAGACTTTATGGGTGTGTTAGAAACAAAGCTGTCGTCTATAGCAGTATCCAAATCGTCTGCTATAGGCAGCTCTTCCTTTTTCTTTTGACCACTATTGCAAGTTCTTAGCCAATCATCGTACTTGATTAGATTGTCTATATTATCATCTTGTTCTTTTGCCATATTTTCACGATCATTCTTTTCAACAGCGTTTGAATACATCGCTTTATAAAACAAAACATATGCTGTTGCCATATTTGGAGATTCACCTGTGAATTCTAACACTGTTTCCTCTTTAAC
 tpg|BK006936.2| 595207 + tpg|BK006936.2| 594647 - INS GCGTTAATGTTGTTTTGATGAACATTAAGCAGGTTACTCATATCAACAGAAGAGTATTCGTAGAATGTATTATTGGATCCTAAAATAATGACAGCAATGTCTACTTGGCAAAGTACTGACAATTCATGAGCCTTTTTAAATAGTCCTGCTTTTCGCTTTATGAAAGTAACTGTACGA
 tpg|BK006945.2| 320872 + tpg|BK006945.2| 321040 - INS GTTCTCTTCCCTGGCGAGTATGATGCGTACGAAGAGGGCAACTCTACAAGCTCTAAGGATATCGATATCGATATATCTCTTACTTTGAAGGATTTGTACATGGGCAAGAAGCTGAAGTTTGATTTAAAGAGACAGGTCATCTGTATAAAGTGCCACGGTTCTGGCTGGAAACCAAAGAGGAAAATTCACGTTACACACGATGTGGAATGTGAATCATGCGCTGGAAAGGGTTCAAAGGAACGTCTGAAG
 tpg|BK006945.2| 754475 + tpg|BK006945.2| 754573 - INS GTACTTTTTGAAACTCTTGCTCTTGAAAAGGTACTGTTATGAGAAGGACGGTTGAAAGGTGTAAAAACTGAACCAGACGCGGCACTGCTTGCTTTTAAATCAATTTGGGAATTTGTTTCTGAATTAGCGCTATATCCTGACGCAGAGGCAATAGCATCTGCCATCTTTGGTGGAATCCTTGATATTGAGGAATTTTTGGACGACGAAGCGGTCACTTCATTAGATGTGACAGCTTTGTTCTTTGTCGCATTACCAAATTCATCCGTAATAAAAGTCGAAAATGGATTTGTCCAAGAACCACCGCTAAATGAACCTTTAAAAAATCTTGGGAGCAACTGTGGTAAAGTATTATCATCTGAGAAGACTGAGCTCTGTAACACAAAATAAAGTAACTGAACATGCCTTAAAAATTTCGAGAATTCCACATCAACCATTTCGTAAATCGATTTAGCTGACTTAAAA
 tpg|BK006945.2| 283644 + tpg|BK006945.2| 283754 - INS CGTCTAACACTGTTGCTTTTTGGATACCAGCAGGAAAAAAAAAAGCCGGAGCTGCAGTAACGAAGAATTGTTGAATGCGTCTAACAAGAAAGGGAGCAATCGATAACAGGGACGTGCGCCGCTAATGTCATTCAGATTATTCACGAGGACTTCTCAACGTCTCCCTCGCCTTAACTGGGTTAGTCCCATCAGGCGATACGCCAAACAACCTCAATACGATGAAGCAGAGTTGTTTGCAGAGAACATTAACCATGGCGCATATAAAGCAAAGAAAAGGCCATCAGACGAGCATTTCCAATGGCCTGAGAAGTCTCCTGATCAGATCACAAAGGAATCTGAACTCCAATGGGAAAGG
 tpg|BK006944.2| 516198 + tpg|BK006944.2| 516220 - INS ATGTACTAGCCTTGTCTGGGTTGTCATCTCTATTCACATGGGGTGGTATCTGTATTTGTCACATTCGTTTCAGAAAGGCATTGGCCGCCCAAGGAAGAGGCTTGGATGAATTGTCTTTCAAGTCTCCTACCGGTGTTTGGGGTTCCTACTGGGGGTTATTTATGGTTATTATTATGTTCATTGCCCAATTCTACGTTGCTGTATTCCCCGTGGGAGATTCTCCAAGTGCGGAAGGTTTCTTCGAAGCTTATC
 tpg|BK006949.2| 911163 + tpg|BK006949.2| 910389 - INS GACTTAAACCCTGATGTACGCTTAATTGGTGTTCAGTCAAAATTGAAGGTCTTGTAAATGCCTTATCACAGCCATCATAGTCACAGAAATATGTCTTTGGCCTATTGCTCGATGAGCTTCTAGTTGATGTTAAACTGTTCAATGATTCTGAACTCTCTGATCGTGATATGGGAATGGTCTCCTGTTTAAGTTCGGCCAGTGGCATTCCTTCATTATTTAGAACCTCTCCTCCCATTTGACAGCGATTTCACCAGTTACTAC
 tpg|BK006944.2| 645848 + tpg|BK006944.2| 646393 - INS GATCCGCTTCCCAGGTTGTACCAGTGAAGCGTGGCGTTAAACTTTGTTCTGATAATACAACTCTTTCTTCTAAAACTGAGAAACGTGAAAATGACGATTGCGATCAAGGCGCTGCCTACTGGAGTTCAGATCTGTTCGGATTCTACACAACACCCACCAACGTAACCGTGGAAATGACAGGTTACTTTTTACCACCAAAAACTGGTACCTACACATTTGGCTTCGCTACTGTGGATGATTCAGCAATTTTATCGGTTGGAGGTAATGTTGCCTTTGAATGTTGTAAACAGGAACAGCCTCCTATCACATCAACGGATT
 tpg|BK006944.2| 142086 + tpg|BK006944.2| 142334 - INS GTTTTAGTGTTGGTAGTGGCTTGGATTTGACCGTCACCAATTTGAGAGACAGCAGCAGCTTTGGTTTTAGTAGTGGCTTGAATGTGACCGTCACCAATTTGGGAGACGGCTGCAGCGGTAGTCTTAGCTGAGGTAGTCTTGGTGGTGGCTTGGATTTGGCCGTCACCAATTTGAGAGACAGCAGCAGCTTTGGTTTTAGTAGTGGCTTGGATTTGACCGTCACCAATTTGAGAAACAGCAGCAGCAGTGGTTTTGGTAGTGGCTTGGATTTGACCGTCACCAATTTGAGAGATAGCAGCGGCTCTCTTAGCCTTGGAG
 tpg|BK006949.2| 283943 + tpg|BK006949.2| 283402 - INS GCAAGGTCTAAAGTACATTTATTTTGCACCATCGTTGGTGCAGGCAGGTCTTTTGAGACTTGATGGGATGTTTGCATATTTGAAGCAGTGATATAATGATTCTTTGAATTTGTTTGATAACTGTCATCCTTTTTTGGGCGTCTTTGGGAAGGTGGAGAAGGTTTCCGTTTGGAATCCATTGATGAGTATAAACTAGATTTGGAAGTATCATAAGAGTACAAGGAAAGAAAGCTAAATCTTTTCTTTGTTGACTCTGCTTCGTTAAGTGATCTTTCTAGATGGTTATTGACGTGTTTTTGTGCTGTAGCTTTCGCGATGTTGCTACTTTTACTACCCTTTTCACTTGTGTCC
 tpg|BK006949.2| 634159 + tpg|BK006949.2| 633625 - INS ACTCTTTTCTTTACTCTTTAGCATTTCAATACCGAACTAAATATCCGTTTTTATAGTTTAGTTGGTTTTGTTTAATTTCTAGAATCCTGTTCGGCGCTTTTGTTAAAAGTAAAAAATGAAAATTCAAACGAAATGAACCTAATCACGTTAGAATTTAAATCTTGGAATATGTTAAATATAAAACAAGAAGAGCAAGCAATACTATTTCTGACTAATTCTCTATACACATAAGAGC
 tpg|BK006949.2| 312473 + tpg|BK006949.2| 312144 - INS GTTAATACAAAGACGGTCAGTGAGTTCACGTTAGACTCTGAAATCCAAACCGTCAAGTTGATTAATGACACAAATTTAATAGTGGCCACCAGGACTACATTAAACGCCATCAACTTATTGCGGGGTCAAGTCATAAATAGTTTTGACTTATATCCGTTTGTTAACGGAGTGTATAAAAA
 tpg|BK006949.2| 197098 + tpg|BK006949.2| 197444 - INS AATTGCTCATTTCGCTGCTTTGTCTGGCATTGAGTTGGTTGCTGTTGAATACGCTGATAATCAAAAATTCCGTCATTCTCGTAAAAGAACGAATCATTAGGCTCTCGTGTAAAGTCGGATGGTAAAAGAGTAAAATTACCATTCATAGGATACACAGCATCGCCAAAGTTTTGAGGGCCACTCGCATAAGTTTCTTGGTAAGGGCCGGAAGAACTGGACTGTTGATACATTGCAAAGTCATCGGAAGAAGGAAAAGGAGGGAACATGTTATTATTG
 tpg|BK006948.2| 278151 + tpg|BK006948.2| 278627 - INS GATGATTGCAATAACGAAAATAGATAGAATTCCACAGCCAAAAGAACGTGAAAAAAAAATTGAAAAAGTTATAAATGATTTGATTGTTCAAGGAATACCAGTAGAGAAAATTGGCGGAGACGTTCAAGTGATCCCGATAAGTGCCAAAACTGGTGAGAAC
 tpg|BK006948.2| 12154 + tpg|BK006948.2| 11586 - INS CTGTTGGGGTCTTTGGAGTATCGTCTCGTGGGCTCGGAGATGTGTATAGAGACAGGAGCTAGAGTGGTGGTTGCGGAAGCACCAGCAGCGATGGCGGCGACACCAGCAGCGATTGAAGTTAATTTGACCATTATATTTGTTTTGTTTTTTAGTGCTGATATGAGCTTAACAGGAAAGAAAGGAATAAAAAAATATTCTCAAAGACATACAGTTGAAGCAGCTCTATTTATACCCATGCCTTCATCAGTCATCACTACTTAAACGATTTGTTAACAGATGCTCATTTATCACTTCACACCTTTCATGTTTCATCTTTCGCACCATCTTCATCATTAAAAATAAGATGCACTTGTTCCTGAACGAGGCATGCATATATCATGAATTTCTTATGCGAAGGTATTGTTCTATGG
 tpg|BK006948.2| 533922 + tpg|BK006948.2| 534204 - INS GAAGAGAATCAACAACAAAGGAATGAGTCGATTTCATATTATACAAATTTCAACCAGCCACGATATTCCACGGACGCCTCTATCAACTCATTCTTGAACATATCTGATAA
 tpg|BK006948.2| 949539 + tpg|BK006948.2| 949330 - INS ATTAAAGATGAAAAAAAAGAGAAAAAAGAAACGGCCAATCCGTTGATCATGATTAAATAAAATATAGGGTTCTGAATTGTTAGGTTTAATCTGCAAATTATTCAGGTCATCGTTGACTTTTTTGCAGGGCACTAAAAACCGCTAACATAGGACGGTATATTGCTGATTTTAGACTTAACTTCTTGGTGTAGTCGTCTCTGAACATGGCATGATACAGCTTTGGTGGGTCACTAGAACAATTTGAATCTTGCTCAGCACGCTCTGTCTTACGTATATATCCAATTTCAGTTGATTCGAAAGACATGAAAGATTATTAATGTGTGCATTACCCGGATTGTCAATAACTCATATAGTTAGTATACTAATTAACTAACTATATAAC
 tpg|BK006943.2| 24368 + tpg|BK006943.2| 23984 - INS GTTCACCTATACATATATAAATTGCAATTGAAAATAGCGTACAGCGTAAGTTAAGTATCCAATGCTCACATATGAAAAGCAAAAGTAAAAAGAAATATACAAGTTTATTATTCATAAATATCGGCATAACTATTTGTTTCGAAAGATCAGTACGTTTATGTTAAATGTGCTCGTTACTTCAACAAGTAAAGTCTTCCTTCCCATGGCTGCAAGGTGCGGGAATCACCATTTGAGTTTGCATAGTTGCCAAAAAACATGGTGTAGGAGGCCTCATTATCAGGAAC
 tpg|BK006943.2| 489233 + tpg|BK006943.2| 488538 - INS GTCTTCATTTCCATGATGGTCTTCAGGCATTACTATTTCCTTAACTTTGATGGACGTGTAAATTTTATGCAAATACCAACGAGGAAAATCTTTTCCATTGTAGCATCCTCGTAAATTGTTAGAGTAGTCATCAAAAGTCATATGGTCTTTAACCTGCGGGTTATGTGAATCGGTATTTAACATGATTATCGAATAACTTAACACAAACACAGAGTCTGCATCAGGCTGTACATGAATGATGTCATCTTCTGTCATTGACTCTGAGCCATTTTTTCCTGCTTTTTTATCCTCTAACTCCACTTTATCATTGCTTTGATCAGCAG
 tpg|BK006943.2| 358890 + tpg|BK006943.2| 358522 - INS ACCTTACACCTTACACAGGTCTAAAAACTTTTCATCATCTTTACTGGCATCTTCCTTTTCAAAAATTTTCTTGAAATGCAAAATCAATTCAACAAATTCATCGTTATTATTCGTATGTTCATAGTCACCTTGGCTCACTAGTTCGTGAAGCTCATCGTAAATGGATAACAAAAGGGTGATGATAGTGCATGCAATGAAAATATCCAAGGGATAATTGAACGTCAGGACGTGGTCCCAAACGATTAGCACATATTTTAAGGGTAATTCTCTTAAAAATAACAACC
