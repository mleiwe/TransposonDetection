NO_ID tpg|BK006942.2| 141108 + tpg|BK006942.2| 141199 - INS
NO_ID tpg|BK006941.2| 467290 + tpg|BK006941.2| 467300 - INS
NO_ID tpg|BK006941.2| 634191 + tpg|BK006941.2| 634308 - INS
NO_ID tpg|BK006941.2| 707252 + tpg|BK006941.2| 706962 - INS
NO_ID tpg|BK006938.2| 1247993 + tpg|BK006938.2| 1248461 - INS
NO_ID tpg|BK006938.2| 221439 + tpg|BK006938.2| 221057 - INS
NO_ID tpg|BK006938.2| 370786 + tpg|BK006938.2| 371454 - INS
NO_ID tpg|BK006938.2| 797664 + tpg|BK006938.2| 798022 - INS
NO_ID tpg|BK006946.2| 917909 + tpg|BK006946.2| 918104 - INS
NO_ID tpg|BK006945.2| 530931 + tpg|BK006945.2| 530751 - INS
NO_ID tpg|BK006945.2| 867286 + tpg|BK006945.2| 867097 - INS
NO_ID tpg|BK006944.2| 310924 + tpg|BK006944.2| 311595 - INS
NO_ID tpg|BK006944.2| 294904 + tpg|BK006944.2| 294351 - INS
NO_ID tpg|BK006949.2| 132924 + tpg|BK006949.2| 133456 - INS
NO_ID tpg|BK006949.2| 838602 + tpg|BK006949.2| 839125 - INS
NO_ID tpg|BK006948.2| 413257 + tpg|BK006948.2| 413040 - INS
NO_ID tpg|BK006943.2| 667739 + tpg|BK006943.2| 667125 - INS
NO_ID tpg|BK006943.2| 53109 + tpg|BK006943.2| 53271 - INS
