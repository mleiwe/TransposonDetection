NO_ID tpg|BK006935.2| 27489 + tpg|BK006935.2| 27084 - INS HAS_CYCLE
NO_ID tpg|BK006935.2| 25652 + tpg|BK006935.2| 25057 - INS HAS_CYCLE
NO_ID tpg|BK006937.2| 152198 + tpg|BK006937.2| 151669 - INS HAS_CYCLE
NO_ID tpg|BK006934.2| 1909 + tpg|BK006934.2| 1805 - INS HAS_CYCLE
NO_ID tpg|BK006941.2| 519207 + tpg|BK006941.2| 518868 - INS HAS_CYCLE
